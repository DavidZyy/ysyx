/* general registers */

`include "./include/defines.v"

module RegisterFile #(ADDR_WIDTH = `RegCnt, DATA_WIDTH = `RegWidth) (
  input clk,
  input [DATA_WIDTH-1:0] wdata,
  input [ADDR_WIDTH-1:0] waddr,
  input wen
);
  reg [DATA_WIDTH-1:0] rf [ADDR_WIDTH-1:0];
  always @(posedge clk) begin
    if (wen) rf[waddr] <= wdata;
  end
endmodule
