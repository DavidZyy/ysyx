`include "defines.v"

/* assemble all cpu moudules into top moudule */
module top(
  input clk,
  input rst,
  input [`InstWidth-1:0] inst
);


endmodule
