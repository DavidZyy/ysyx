// soc(system on chip)

`include "./include/defines.v"

module top	(
        input	clk,
        input	sysclk_n,
        /* verilator lint_off SYNCASYNCNET */
        input 	rst,
		/* verilator lint_off UNUSEDSIGNAL */
        // input	btn_clk,
        input   PS2_clk,
        input   PS2_Data,
        input   [`Vec(8)]   swt,

        // output  [`Vec(`ImmWidth)] pc_WB,
        // output  [`Vec(`ImmWidth)] pc_IF,
        // output  flush_WB,
        output	[7:0] leds,
        output  SEGCLK,
        output  SEGCLR,
        output  SEGDT,
        output  SEGEN,
        output  [3:0]   vga_r,
        output  [3:0]   vga_g,
        output  [3:0]   vga_b,
        output  vga_hs,
        output  vga_vs
);

    /* verilator lint_off UNUSEDSIGNAL */
    wire [`Vec(`ImmWidth)] pc_WB;
    wire [`Vec(`ImmWidth)] pc_IF;
    wire flush_WB;
    wire [`Vec(`InstWidth)]	inst;

    wire    clk200m;
    reg [`Vec(`ClkDivWidth)]  clkdiv;

    IBUFDS  inst_clk(
                .I(clk),
                .IB(sysclk_n),

                .O(clk200m)
            );

    /* seg no display, to see rst signal */
    always@(posedge clk200m or posedge rst) begin
      if(rst) begin
    	clkdiv <= 0;
      end
      else begin
        clkdiv <= clkdiv+1;
      end
    end
    	
    // wire clk100m = clkdiv[0];
    // wire clk50m  = clkdiv[1];
    // wire clk25m  = clkdiv[2];
    // wire clk12m  = clkdiv[3];

    wire clk100m;
    wire clk50m ;
    wire clk25m ;

    divider #(2) div1(clk200m, rst, clk100m);
    divider #(4) div2(clk200m, rst, clk50m );
    divider #(8) div3(clk200m, rst, clk25m );

    wire sig_rd_kb;
    wire [`Vec(`SegWidth)]  seg_wdata;

    wire [`Vec(`KbWidth)]	kb_rdata;
    wire kb_ready;
    wire overflow;

    wire [`Vec(`LedWidth)]	led_wdata;

    wire [`Vec(8)]	swt_rdata;
    cpu u_cpu (
            //ports
            .cpu_clk        	( clk25m			), /* for simulation on varilator */
            .clkdiv             ( clkdiv            ),
            /* 10 can run on sword */
            // .cpu_clk        	( clkdiv[10]		),
            // .clk        		( btn_clk			),
            /* use switch as reset? */
            .rst        		( rst        		),
            .kb_rdata     		( kb_rdata     		),
            .kb_ready    		( kb_ready    		),
            .swt_rdata          ( swt_rdata         ),

            .inst           	( inst 				),
            .pc_IF				( pc_IF				),
            .flush_WB			( flush_WB			),
            .pc_WB				( pc_WB				),
            .sig_rd_kb			( sig_rd_kb			),
            .seg_wdata			( seg_wdata			),
            .led_wdata          ( led_wdata         )
        );

    // always@(posedge clk200m) begin
    // 	$display("%x", pc_WB);
    // end

//     assign leds[7] = btn_clk;
//     /* rst always true */
//     assign leds[6] = rst;
//     assign leds[5] = flush_WB;
//     assign leds[4] = clk200m;
// 
//     assign leds[3:0] = pc_IF[3:0];


    swt u_swt (
    	//ports
    	.swt       		( swt       		),

    	.swt_rdata 		( swt_rdata 		)
    );


	assign leds [6:0] = led_wdata[6:0];
	// assign leds [5:0] = led_wdata[5:0];
	// assign leds [4:0] = led_wdata[4:0];
    // assign leds[5] = swt_rdata[5];
    // assign leds[6] = swt[6];
    assign leds[7] = rst;
//     led u_led (
//     	//ports
//     	.led_wdata 		( led_wdata 		),
//     	// .led_wdata 		( seg_wdata[7:0] ),
// 
//     	.led_out   		( leds           )
//     );

    wire [`Vec(`ImmWidth)] led_ext = `ZEXT(led_wdata, 8);

    // seg_wdata shift left to display the signal
    // reg [`Vec(`SegWidth)] seg_wdata2;
    // always @(*) begin
    //     if(rst)
    //         seg_wdata2 = 0;
    //     else
    //         seg_wdata2 = {seg_wdata2[23:0], seg_wdata[7:0]};
    // end

    seg u_seg (
            //ports
            .clkdiv   		( clkdiv   		),
            // .num    		( seg_wdata2	),
            .num    		( seg_wdata	    ),

            .s_clk  		( SEGCLK		),
            .s_clrn 		( SEGCLR		),
            .sout   		( SEGDT			),
            .EN     		( SEGEN		    )
        );

    ps2_kbd u_ps2_kbd (
                //ports
                /* clk200m may be too quickly? */
                // .kb_clk      	( clk25m       ),
                .kb_clk      	( clk200m       ),
                .clrn     		( rst			),
                .ps2_clk  		( PS2_clk  		),
                .ps2_data 		( PS2_Data 		),
                .rdn      		( sig_rd_kb     ),

                .data     		( kb_rdata     	),
                .ready    		( kb_ready    	),
                .overflow       ( overflow      )
            );

    wire [8:0]	row;
    wire [9:0]	col;
    wire rdn;

    // wire [3:0]	R;
    // wire [3:0]	G;
    // wire [3:0]	B;
    // wire HS;
    // wire VS;

    VGA u_VGA(
    	//ports
    	.clk 		( clk25m    ),
    	.rst 		( rst 		),
    	.din 		( 12'b0     ),

    	.row 		( row 		),
    	.col 		( col 		),
    	.rdn 		( rdn 		),
    	.R   		( vga_r   	),
    	.G   		( vga_g   	),
    	.B   		( vga_b   	),
    	.HS  		( vga_hs    ),
    	.VS  		( vga_vs    )
    );

endmodule //top
