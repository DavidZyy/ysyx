/* verilator lint_off DECLFILENAME */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off UNDRIVEN */
/* verilator lint_off UNOPTFLAT */
/* verilator lint_off WIDTHEXPAND */
module IDU(
  input         from_IFU_valid,
  input  [31:0] from_IFU_bits_inst,
  input  [31:0] from_IFU_bits_pc,
  output        to_ISU_valid,
  output [31:0] to_ISU_bits_imm,
  output [31:0] to_ISU_bits_pc,
  output [4:0]  to_ISU_bits_rs1,
  output [4:0]  to_ISU_bits_rs2,
  output [4:0]  to_ISU_bits_rd,
  output        to_ISU_bits_ctrl_sig_reg_wen,
  output [2:0]  to_ISU_bits_ctrl_sig_fu_op,
  output        to_ISU_bits_ctrl_sig_mem_wen,
  output        to_ISU_bits_ctrl_sig_is_ebreak,
  output        to_ISU_bits_ctrl_sig_not_impl,
  output [1:0]  to_ISU_bits_ctrl_sig_src1_op,
  output [1:0]  to_ISU_bits_ctrl_sig_src2_op,
  output [3:0]  to_ISU_bits_ctrl_sig_alu_op,
  output [3:0]  to_ISU_bits_ctrl_sig_lsu_op,
  output [3:0]  to_ISU_bits_ctrl_sig_bru_op,
  output [2:0]  to_ISU_bits_ctrl_sig_csr_op,
  output [3:0]  to_ISU_bits_ctrl_sig_mdu_op
);
  wire [19:0] _imm_i_T_2 = from_IFU_bits_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_i = {_imm_i_T_2,from_IFU_bits_inst[31:20]}; // @[Cat.scala 33:92]
  wire [31:0] imm_s = {_imm_i_T_2,from_IFU_bits_inst[31:25],from_IFU_bits_inst[11:7]}; // @[Cat.scala 33:92]
  wire [31:0] imm_b = {_imm_i_T_2,from_IFU_bits_inst[7],from_IFU_bits_inst[30:25],from_IFU_bits_inst[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] imm_u = {from_IFU_bits_inst[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [11:0] _imm_j_T_2 = from_IFU_bits_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 77:12]
  wire [32:0] imm_j = {_imm_j_T_2,from_IFU_bits_inst[31],from_IFU_bits_inst[19:12],from_IFU_bits_inst[20],
    from_IFU_bits_inst[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] decode_info_invInputs = ~from_IFU_bits_inst; // @[pla.scala 78:21]
  wire  decode_info_andMatrixInput_0 = from_IFU_bits_inst[0]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_1 = from_IFU_bits_inst[1]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_2 = decode_info_invInputs[2]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_3 = decode_info_invInputs[3]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_4 = decode_info_invInputs[4]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_5 = decode_info_invInputs[5]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_6 = decode_info_invInputs[6]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_7 = decode_info_invInputs[13]; // @[pla.scala 91:29]
  wire [7:0] _decode_info_T = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_1 = &_decode_info_T; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_6_1 = decode_info_invInputs[12]; // @[pla.scala 91:29]
  wire [7:0] _decode_info_T_2 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_3 = &_decode_info_T_2; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_7_2 = decode_info_invInputs[14]; // @[pla.scala 91:29]
  wire [7:0] _decode_info_T_4 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_5 = &_decode_info_T_4; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_6 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_7 = &_decode_info_T_6; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_8 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_9 = &_decode_info_T_8; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_10 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_6,decode_info_andMatrixInput_7
    ,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_11 = &_decode_info_T_10; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_4_6 = from_IFU_bits_inst[4]; // @[pla.scala 90:45]
  wire [7:0] _decode_info_T_12 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1}; // @[Cat.scala 33:92]
  wire  _decode_info_T_13 = &_decode_info_T_12; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_2_7 = from_IFU_bits_inst[2]; // @[pla.scala 90:45]
  wire [5:0] _decode_info_T_14 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_info_T_15 = &_decode_info_T_14; // @[pla.scala 98:74]
  wire [6:0] _decode_info_T_16 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_info_T_17 = &_decode_info_T_16; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_5_9 = from_IFU_bits_inst[5]; // @[pla.scala 90:45]
  wire [8:0] _decode_info_T_18 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_19 = &_decode_info_T_18; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_20 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_21 = &_decode_info_T_20; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_22 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_23 = &_decode_info_T_22; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_10 = decode_info_invInputs[25]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_11 = decode_info_invInputs[26]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_12 = decode_info_invInputs[27]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_13 = decode_info_invInputs[28]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_14 = decode_info_invInputs[29]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_15 = decode_info_invInputs[31]; // @[pla.scala 91:29]
  wire [7:0] decode_info_lo_12 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2,
    decode_info_andMatrixInput_10,decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,
    decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_24 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_12}; // @[Cat.scala 33:92]
  wire  _decode_info_T_25 = &_decode_info_T_24; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_11_1 = decode_info_invInputs[30]; // @[pla.scala 91:29]
  wire [5:0] decode_info_lo_13 = {decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,
    decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,
    decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [12:0] _decode_info_T_26 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_lo_13}; // @[Cat.scala 33:92]
  wire  _decode_info_T_27 = &_decode_info_T_26; // @[pla.scala 98:74]
  wire [6:0] decode_info_lo_14 = {decode_info_andMatrixInput_10,decode_info_andMatrixInput_11,
    decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,
    decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_T_28 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_lo_14}; // @[Cat.scala 33:92]
  wire  _decode_info_T_29 = &_decode_info_T_28; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_15 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_30 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_15}; // @[Cat.scala 33:92]
  wire  _decode_info_T_31 = &_decode_info_T_30; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_6_15 = from_IFU_bits_inst[6]; // @[pla.scala 90:45]
  wire [7:0] _decode_info_T_32 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_33 = &_decode_info_T_32; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_34 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_35 = &_decode_info_T_34; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_36 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_3
    ,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_37 = &_decode_info_T_36; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_38 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_39 = &_decode_info_T_38; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_3_20 = from_IFU_bits_inst[3]; // @[pla.scala 90:45]
  wire [6:0] _decode_info_T_40 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3_20,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15}; // @[Cat.scala 33:92]
  wire  _decode_info_T_41 = &_decode_info_T_40; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_7_18 = decode_info_invInputs[7]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_8_10 = decode_info_invInputs[8]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_9_5 = decode_info_invInputs[9]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_10_4 = decode_info_invInputs[10]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_11_4 = decode_info_invInputs[11]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_15_2 = decode_info_invInputs[15]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_16 = decode_info_invInputs[16]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_17 = decode_info_invInputs[17]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_18 = decode_info_invInputs[18]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_19 = decode_info_invInputs[19]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_20 = decode_info_invInputs[21]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_21 = decode_info_invInputs[22]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_22 = decode_info_invInputs[23]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_23 = decode_info_invInputs[24]; // @[pla.scala 91:29]
  wire [14:0] decode_info_lo_21 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,decode_info_andMatrixInput_20,
    decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_andMatrixInput_23,decode_info_lo_14}; // @[Cat.scala 33:92]
  wire [7:0] decode_info_hi_lo_20 = {decode_info_andMatrixInput_8_10,decode_info_andMatrixInput_9_5,
    decode_info_andMatrixInput_10_4,decode_info_andMatrixInput_11_4,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_15_2}; // @[Cat.scala 33:92]
  wire [30:0] _decode_info_T_42 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_21}; // @[Cat.scala 33:92]
  wire  _decode_info_T_43 = &_decode_info_T_42; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_20_1 = decode_info_invInputs[20]; // @[pla.scala 91:29]
  wire [7:0] decode_info_lo_lo_19 = {decode_info_andMatrixInput_23,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] decode_info_lo_22 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,decode_info_andMatrixInput_20_1,
    decode_info_andMatrixInput_20,decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_lo_lo_19}; // @[Cat.scala 33:92]
  wire [31:0] _decode_info_T_44 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_22}; // @[Cat.scala 33:92]
  wire  _decode_info_T_45 = &_decode_info_T_44; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_6_22 = from_IFU_bits_inst[12]; // @[pla.scala 90:45]
  wire [8:0] _decode_info_T_46 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_47 = &_decode_info_T_46; // @[pla.scala 98:74]
  wire [6:0] decode_info_lo_24 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_11,
    decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,
    decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_T_48 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_24}; // @[Cat.scala 33:92]
  wire  _decode_info_T_49 = &_decode_info_T_48; // @[pla.scala 98:74]
  wire [14:0] _decode_info_T_50 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_24}; // @[Cat.scala 33:92]
  wire  _decode_info_T_51 = &_decode_info_T_50; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_52 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_53 = &_decode_info_T_52; // @[pla.scala 98:74]
  wire [15:0] _decode_info_T_54 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_15}; // @[Cat.scala 33:92]
  wire  _decode_info_T_55 = &_decode_info_T_54; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_56 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_57 = &_decode_info_T_56; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_58 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,
    decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_59 = &_decode_info_T_58; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_60 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_61 = &_decode_info_T_60; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_8_20 = from_IFU_bits_inst[13]; // @[pla.scala 90:45]
  wire [9:0] _decode_info_T_62 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6
    ,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_63 = &_decode_info_T_62; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_64 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_8_20}; // @[Cat.scala 33:92]
  wire  _decode_info_T_65 = &_decode_info_T_64; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_66 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_67 = &_decode_info_T_66; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_68 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_20,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_69 = &_decode_info_T_68; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_35 = {decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_70 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_8_20,decode_info_lo_35}; // @[Cat.scala 33:92]
  wire  _decode_info_T_71 = &_decode_info_T_70; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_72 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_20,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_73 = &_decode_info_T_72; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_74 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_8_20}; // @[Cat.scala 33:92]
  wire  _decode_info_T_75 = &_decode_info_T_74; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_38 = {decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_76 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_38}; // @[Cat.scala 33:92]
  wire  _decode_info_T_77 = &_decode_info_T_76; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_8_27 = from_IFU_bits_inst[14]; // @[pla.scala 90:45]
  wire [8:0] _decode_info_T_78 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6
    ,decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_79 = &_decode_info_T_78; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_80 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_81 = &_decode_info_T_80; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_41 = {decode_info_andMatrixInput_8_27,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_82 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_41}; // @[Cat.scala 33:92]
  wire  _decode_info_T_83 = &_decode_info_T_82; // @[pla.scala 98:74]
  wire [15:0] _decode_info_T_84 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_7,decode_info_lo_41}; // @[Cat.scala 33:92]
  wire  _decode_info_T_85 = &_decode_info_T_84; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_86 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_87 = &_decode_info_T_86; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_88 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_89 = &_decode_info_T_88; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_90 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6
    ,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_91 = &_decode_info_T_90; // @[pla.scala 98:74]
  wire [6:0] decode_info_lo_46 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [14:0] _decode_info_T_92 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_46}; // @[Cat.scala 33:92]
  wire  _decode_info_T_93 = &_decode_info_T_92; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_47 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_94 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_47}; // @[Cat.scala 33:92]
  wire  _decode_info_T_95 = &_decode_info_T_94; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_48 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_10,decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,
    decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_96 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_48}; // @[Cat.scala 33:92]
  wire  _decode_info_T_97 = &_decode_info_T_96; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_98 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,
    decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_99 = &_decode_info_T_98; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_100 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_101 = &_decode_info_T_100; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_102 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_103 = &_decode_info_T_102; // @[pla.scala 98:74]
  wire [15:0] decode_info_lo_52 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,from_IFU_bits_inst[20],decode_info_andMatrixInput_20,
    decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_lo_lo_19}; // @[Cat.scala 33:92]
  wire [31:0] _decode_info_T_104 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_52}; // @[Cat.scala 33:92]
  wire  _decode_info_T_105 = &_decode_info_T_104; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_7_50 = from_IFU_bits_inst[25]; // @[pla.scala 90:45]
  wire [6:0] decode_info_lo_53 = {decode_info_andMatrixInput_7_50,decode_info_andMatrixInput_11,
    decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,
    decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_T_106 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_lo_53}; // @[Cat.scala 33:92]
  wire  _decode_info_T_107 = &_decode_info_T_106; // @[pla.scala 98:74]
  wire [14:0] _decode_info_T_108 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_53}; // @[Cat.scala 33:92]
  wire  _decode_info_T_109 = &_decode_info_T_108; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_55 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_110 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_55}; // @[Cat.scala 33:92]
  wire  _decode_info_T_111 = &_decode_info_T_110; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_56 = {decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_112 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_56}; // @[Cat.scala 33:92]
  wire  _decode_info_T_113 = &_decode_info_T_112; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_57 = {decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [16:0] _decode_info_T_114 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_8_20,decode_info_lo_57}; // @[Cat.scala 33:92]
  wire  _decode_info_T_115 = &_decode_info_T_114; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_58 = {decode_info_andMatrixInput_8_27,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_116 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_58}; // @[Cat.scala 33:92]
  wire  _decode_info_T_117 = &_decode_info_T_116; // @[pla.scala 98:74]
  wire [15:0] _decode_info_T_118 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_7,decode_info_lo_58}; // @[Cat.scala 33:92]
  wire  _decode_info_T_119 = &_decode_info_T_118; // @[pla.scala 98:74]
  wire [16:0] _decode_info_T_120 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_8_20,decode_info_lo_58}; // @[Cat.scala 33:92]
  wire  _decode_info_T_121 = &_decode_info_T_120; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_21_3 = from_IFU_bits_inst[21]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_28_3 = from_IFU_bits_inst[28]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_29_3 = from_IFU_bits_inst[29]; // @[pla.scala 90:45]
  wire [7:0] decode_info_lo_lo_58 = {decode_info_andMatrixInput_23,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_28_3,
    decode_info_andMatrixInput_29_3,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] decode_info_lo_61 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,decode_info_andMatrixInput_20_1,
    decode_info_andMatrixInput_21_3,decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_lo_lo_58}; // @[Cat.scala 33:92]
  wire [31:0] _decode_info_T_122 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_61}; // @[Cat.scala 33:92]
  wire  _decode_info_T_123 = &_decode_info_T_122; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_15_19 = from_IFU_bits_inst[30]; // @[pla.scala 90:45]
  wire [7:0] decode_info_lo_62 = {decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15_19,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [16:0] _decode_info_T_124 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_7,decode_info_lo_62}; // @[Cat.scala 33:92]
  wire  _decode_info_T_125 = &_decode_info_T_124; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_63 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15_19,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_126 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_63}; // @[Cat.scala 33:92]
  wire  _decode_info_T_127 = &_decode_info_T_126; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_64 = {decode_info_andMatrixInput_8_27,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15_19,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [16:0] _decode_info_T_128 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_7,decode_info_lo_64}; // @[Cat.scala 33:92]
  wire  _decode_info_T_129 = &_decode_info_T_128; // @[pla.scala 98:74]
  wire  _decode_info_orMatrixOutputs_T = |_decode_info_T_109; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_1 = {_decode_info_T_111,_decode_info_T_113}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_2 = |_decode_info_orMatrixOutputs_T_1; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_3 = {_decode_info_T_115,_decode_info_T_117,_decode_info_T_119}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_4 = |_decode_info_orMatrixOutputs_T_3; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_5 = |_decode_info_T_121; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_6 = {_decode_info_T_45,_decode_info_T_61}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_7 = |_decode_info_orMatrixOutputs_T_6; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_8 = {_decode_info_T_61,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_9 = |_decode_info_orMatrixOutputs_T_8; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_10 = |_decode_info_T_73; // @[pla.scala 114:39]
  wire [8:0] decode_info_orMatrixOutputs_lo = {_decode_info_T_43,_decode_info_T_49,_decode_info_T_59,_decode_info_T_65,
    _decode_info_T_73,_decode_info_T_87,_decode_info_T_93,_decode_info_T_97,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [17:0] _decode_info_orMatrixOutputs_T_11 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_11,
    _decode_info_T_15,_decode_info_T_25,_decode_info_T_27,_decode_info_T_37,_decode_info_T_41,
    decode_info_orMatrixOutputs_lo}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_12 = |_decode_info_orMatrixOutputs_T_11; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_13 = |_decode_info_T_105; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_14 = {_decode_info_T_19,_decode_info_T_23}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_15 = |_decode_info_orMatrixOutputs_T_14; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_1 = {_decode_info_T_41,_decode_info_T_49,_decode_info_T_61,_decode_info_T_65
    ,_decode_info_T_73,_decode_info_T_93,_decode_info_T_97}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_orMatrixOutputs_T_16 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_7,_decode_info_T_15,
    _decode_info_T_25,_decode_info_T_27,_decode_info_T_39,decode_info_orMatrixOutputs_lo_1}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_17 = |_decode_info_orMatrixOutputs_T_16; // @[pla.scala 114:39]
  wire [4:0] decode_info_orMatrixOutputs_lo_2 = {_decode_info_T_41,_decode_info_T_51,_decode_info_T_65,_decode_info_T_87
    ,_decode_info_T_93}; // @[Cat.scala 33:92]
  wire [10:0] _decode_info_orMatrixOutputs_T_18 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_15,
    _decode_info_T_21,_decode_info_T_37,decode_info_orMatrixOutputs_lo_2}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_19 = |_decode_info_orMatrixOutputs_T_18; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_3 = {_decode_info_T_37,_decode_info_T_41,_decode_info_T_49,_decode_info_T_65
    ,_decode_info_T_87,_decode_info_T_93,_decode_info_T_97}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_orMatrixOutputs_T_20 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_15,
    _decode_info_T_21,_decode_info_T_25,_decode_info_T_27,decode_info_orMatrixOutputs_lo_3}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_21 = |_decode_info_orMatrixOutputs_T_20; // @[pla.scala 114:39]
  wire [3:0] _decode_info_orMatrixOutputs_T_22 = {_decode_info_T_17,_decode_info_T_33,_decode_info_T_41,
    _decode_info_T_87}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_23 = |_decode_info_orMatrixOutputs_T_22; // @[pla.scala 114:39]
  wire [4:0] decode_info_orMatrixOutputs_lo_5 = {_decode_info_T_39,_decode_info_T_49,_decode_info_T_65,_decode_info_T_93
    ,_decode_info_T_97}; // @[Cat.scala 33:92]
  wire [10:0] _decode_info_orMatrixOutputs_T_24 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_11,
    _decode_info_T_25,_decode_info_T_27,decode_info_orMatrixOutputs_lo_5}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_25 = |_decode_info_orMatrixOutputs_T_24; // @[pla.scala 114:39]
  wire [5:0] decode_info_orMatrixOutputs_lo_6 = {_decode_info_T_41,_decode_info_T_75,_decode_info_T_77,_decode_info_T_85
    ,_decode_info_T_87,_decode_info_T_95}; // @[Cat.scala 33:92]
  wire [12:0] _decode_info_orMatrixOutputs_T_26 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_15,
    _decode_info_T_21,_decode_info_T_31,_decode_info_T_37,decode_info_orMatrixOutputs_lo_6}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_27 = |_decode_info_orMatrixOutputs_T_26; // @[pla.scala 114:39]
  wire [6:0] _decode_info_orMatrixOutputs_T_28 = {_decode_info_T_67,_decode_info_T_71,_decode_info_T_75,
    _decode_info_T_77,_decode_info_T_125,_decode_info_T_127,_decode_info_T_129}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_29 = |_decode_info_orMatrixOutputs_T_28; // @[pla.scala 114:39]
  wire [3:0] _decode_info_orMatrixOutputs_T_30 = {_decode_info_T_67,_decode_info_T_71,_decode_info_T_81,
    _decode_info_T_83}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_31 = |_decode_info_orMatrixOutputs_T_30; // @[pla.scala 114:39]
  wire [3:0] _decode_info_orMatrixOutputs_T_32 = {_decode_info_T_51,_decode_info_T_55,_decode_info_T_93,
    _decode_info_T_97}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_33 = |_decode_info_orMatrixOutputs_T_32; // @[pla.scala 114:39]
  wire [5:0] decode_info_orMatrixOutputs_lo_10 = {_decode_info_T_59,_decode_info_T_65,_decode_info_T_73,
    _decode_info_T_87,_decode_info_T_93,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [11:0] _decode_info_orMatrixOutputs_T_34 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_7,_decode_info_T_37,
    _decode_info_T_41,_decode_info_T_51,decode_info_orMatrixOutputs_lo_10}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_35 = |_decode_info_orMatrixOutputs_T_34; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_11 = {_decode_info_T_49,_decode_info_T_61,_decode_info_T_65,
    _decode_info_T_73,_decode_info_T_93,_decode_info_T_97,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [14:0] _decode_info_orMatrixOutputs_T_36 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_7,_decode_info_T_15,
    _decode_info_T_25,_decode_info_T_27,_decode_info_T_39,_decode_info_T_41,decode_info_orMatrixOutputs_lo_11}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_37 = |_decode_info_orMatrixOutputs_T_36; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_12 = {_decode_info_T_59,_decode_info_T_65,_decode_info_T_73,
    _decode_info_T_87,_decode_info_T_93,_decode_info_T_97,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [14:0] _decode_info_orMatrixOutputs_T_38 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_11,
    _decode_info_T_25,_decode_info_T_27,_decode_info_T_37,_decode_info_T_49,decode_info_orMatrixOutputs_lo_12}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_39 = |_decode_info_orMatrixOutputs_T_38; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_40 = {_decode_info_T_35,_decode_info_T_41,_decode_info_T_89}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_41 = |_decode_info_orMatrixOutputs_T_40; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_42 = {_decode_info_T_37,_decode_info_T_99,_decode_info_T_101}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_43 = |_decode_info_orMatrixOutputs_T_42; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_44 = {_decode_info_T_57,_decode_info_T_89}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_45 = |_decode_info_orMatrixOutputs_T_44; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_46 = |_decode_info_T_103; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_47 = {_decode_info_T_9,_decode_info_T_53,_decode_info_T_91}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_48 = |_decode_info_orMatrixOutputs_T_47; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_49 = {_decode_info_T_23,_decode_info_T_47,_decode_info_T_63}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_50 = |_decode_info_orMatrixOutputs_T_49; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_51 = {_decode_info_T_23,_decode_info_T_79}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_52 = |_decode_info_orMatrixOutputs_T_51; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_53 = |_decode_info_T_69; // @[pla.scala 114:39]
  wire [14:0] _decode_info_orMatrixOutputs_T_54 = {_decode_info_T_13,_decode_info_T_15,_decode_info_T_25,
    _decode_info_T_29,_decode_info_T_37,_decode_info_T_41,_decode_info_T_43,_decode_info_T_51,
    decode_info_orMatrixOutputs_lo_12}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_55 = |_decode_info_orMatrixOutputs_T_54; // @[pla.scala 114:39]
  wire [4:0] _decode_info_orMatrixOutputs_T_56 = {_decode_info_T_33,_decode_info_T_37,_decode_info_T_41,
    _decode_info_T_87,_decode_info_T_107}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_57 = |_decode_info_orMatrixOutputs_T_56; // @[pla.scala 114:39]
  wire [6:0] _decode_info_orMatrixOutputs_T_58 = {_decode_info_T_1,_decode_info_T_5,_decode_info_T_11,_decode_info_T_43,
    _decode_info_T_61,_decode_info_T_73,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_59 = |_decode_info_orMatrixOutputs_T_58; // @[pla.scala 114:39]
  wire [7:0] decode_info_orMatrixOutputs_lo_lo_10 = {_decode_info_orMatrixOutputs_T_12,_decode_info_orMatrixOutputs_T_10
    ,_decode_info_orMatrixOutputs_T_9,_decode_info_orMatrixOutputs_T_7,_decode_info_orMatrixOutputs_T_5,
    _decode_info_orMatrixOutputs_T_4,_decode_info_orMatrixOutputs_T_2,_decode_info_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decode_info_orMatrixOutputs_hi_lo_12 = {_decode_info_orMatrixOutputs_T_43,_decode_info_orMatrixOutputs_T_41
    ,_decode_info_orMatrixOutputs_T_39,_decode_info_orMatrixOutputs_T_37,_decode_info_orMatrixOutputs_T_35,
    _decode_info_orMatrixOutputs_T_33,_decode_info_orMatrixOutputs_T_31,_decode_info_orMatrixOutputs_T_29}; // @[Cat.scala 33:92]
  wire [16:0] decode_info_orMatrixOutputs_hi_21 = {_decode_info_orMatrixOutputs_T_59,_decode_info_orMatrixOutputs_T_57,
    _decode_info_orMatrixOutputs_T_55,_decode_info_orMatrixOutputs_T_53,_decode_info_orMatrixOutputs_T_52,
    _decode_info_orMatrixOutputs_T_50,_decode_info_orMatrixOutputs_T_48,_decode_info_orMatrixOutputs_T_46,
    _decode_info_orMatrixOutputs_T_45,decode_info_orMatrixOutputs_hi_lo_12}; // @[Cat.scala 33:92]
  wire [32:0] decode_info_orMatrixOutputs = {decode_info_orMatrixOutputs_hi_21,_decode_info_orMatrixOutputs_T_27,
    _decode_info_orMatrixOutputs_T_25,_decode_info_orMatrixOutputs_T_23,_decode_info_orMatrixOutputs_T_21,
    _decode_info_orMatrixOutputs_T_19,_decode_info_orMatrixOutputs_T_17,_decode_info_orMatrixOutputs_T_15,
    _decode_info_orMatrixOutputs_T_13,decode_info_orMatrixOutputs_lo_lo_10}; // @[Cat.scala 33:92]
  wire  _decode_info_invMatrixOutputs_T_8 = ~decode_info_orMatrixOutputs[7]; // @[pla.scala 123:40]
  wire  _decode_info_invMatrixOutputs_T_22 = ~decode_info_orMatrixOutputs[20]; // @[pla.scala 123:40]
  wire  _decode_info_invMatrixOutputs_T_24 = ~decode_info_orMatrixOutputs[21]; // @[pla.scala 123:40]
  wire [7:0] decode_info_invMatrixOutputs_lo_lo = {_decode_info_invMatrixOutputs_T_8,decode_info_orMatrixOutputs[6],
    decode_info_orMatrixOutputs[5],decode_info_orMatrixOutputs[4],decode_info_orMatrixOutputs[3],
    decode_info_orMatrixOutputs[2],decode_info_orMatrixOutputs[1],decode_info_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] decode_info_invMatrixOutputs_hi_lo = {decode_info_orMatrixOutputs[23],decode_info_orMatrixOutputs[22],
    _decode_info_invMatrixOutputs_T_24,_decode_info_invMatrixOutputs_T_22,decode_info_orMatrixOutputs[19],
    decode_info_orMatrixOutputs[18],decode_info_orMatrixOutputs[17],decode_info_orMatrixOutputs[16]}; // @[Cat.scala 33:92]
  wire [16:0] decode_info_invMatrixOutputs_hi = {decode_info_orMatrixOutputs[32],decode_info_orMatrixOutputs[31],
    decode_info_orMatrixOutputs[30],decode_info_orMatrixOutputs[29],decode_info_orMatrixOutputs[28],
    decode_info_orMatrixOutputs[27],decode_info_orMatrixOutputs[26],decode_info_orMatrixOutputs[25],
    decode_info_orMatrixOutputs[24],decode_info_invMatrixOutputs_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] decode_info_invMatrixOutputs = {decode_info_invMatrixOutputs_hi,decode_info_orMatrixOutputs[15],
    decode_info_orMatrixOutputs[14],decode_info_orMatrixOutputs[13],decode_info_orMatrixOutputs[12],
    decode_info_orMatrixOutputs[11],decode_info_orMatrixOutputs[10],decode_info_orMatrixOutputs[9],
    decode_info_orMatrixOutputs[8],decode_info_invMatrixOutputs_lo_lo}; // @[Cat.scala 33:92]
  wire [2:0] inst_type = decode_info_invMatrixOutputs[21:19]; // @[IDU.scala 111:36]
  wire [31:0] _to_ISU_bits_imm_T_1 = 3'h1 == inst_type ? imm_i : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_imm_T_3 = 3'h2 == inst_type ? imm_s : _to_ISU_bits_imm_T_1; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_imm_T_5 = 3'h3 == inst_type ? imm_b : _to_ISU_bits_imm_T_3; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_imm_T_7 = 3'h4 == inst_type ? imm_u : _to_ISU_bits_imm_T_5; // @[Mux.scala 81:58]
  wire [32:0] _to_ISU_bits_imm_T_9 = 3'h5 == inst_type ? imm_j : {{1'd0}, _to_ISU_bits_imm_T_7}; // @[Mux.scala 81:58]
  assign to_ISU_valid = from_IFU_valid; // @[IDU.scala 17:20]
  assign to_ISU_bits_imm = _to_ISU_bits_imm_T_9[31:0]; // @[IDU.scala 112:21]
  assign to_ISU_bits_pc = from_IFU_bits_pc; // @[IDU.scala 122:21]
  assign to_ISU_bits_rs1 = from_IFU_bits_inst[19:15]; // @[IDU.scala 119:42]
  assign to_ISU_bits_rs2 = from_IFU_bits_inst[24:20]; // @[IDU.scala 120:42]
  assign to_ISU_bits_rd = from_IFU_bits_inst[11:7]; // @[IDU.scala 121:42]
  assign to_ISU_bits_ctrl_sig_reg_wen = decode_info_invMatrixOutputs[10]; // @[IDU.scala 130:50]
  assign to_ISU_bits_ctrl_sig_fu_op = decode_info_invMatrixOutputs[32:30]; // @[IDU.scala 136:50]
  assign to_ISU_bits_ctrl_sig_mem_wen = decode_info_invMatrixOutputs[9]; // @[IDU.scala 129:50]
  assign to_ISU_bits_ctrl_sig_is_ebreak = decode_info_invMatrixOutputs[8]; // @[IDU.scala 128:50]
  assign to_ISU_bits_ctrl_sig_not_impl = decode_info_invMatrixOutputs[7]; // @[IDU.scala 127:50]
  assign to_ISU_bits_ctrl_sig_src1_op = decode_info_invMatrixOutputs[14:13]; // @[IDU.scala 132:50]
  assign to_ISU_bits_ctrl_sig_src2_op = decode_info_invMatrixOutputs[12:11]; // @[IDU.scala 131:50]
  assign to_ISU_bits_ctrl_sig_alu_op = decode_info_invMatrixOutputs[18:15]; // @[IDU.scala 133:50]
  assign to_ISU_bits_ctrl_sig_lsu_op = decode_info_invMatrixOutputs[29:26]; // @[IDU.scala 135:50]
  assign to_ISU_bits_ctrl_sig_bru_op = decode_info_invMatrixOutputs[25:22]; // @[IDU.scala 134:50]
  assign to_ISU_bits_ctrl_sig_csr_op = decode_info_invMatrixOutputs[6:4]; // @[IDU.scala 126:50]
  assign to_ISU_bits_ctrl_sig_mdu_op = decode_info_invMatrixOutputs[3:0]; // @[IDU.scala 125:50]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_in_rs1,
  input  [4:0]  io_in_rs2,
  input  [4:0]  io_in_rd,
  input  [31:0] io_in_wdata,
  input         io_in_reg_wen,
  output [31:0] io_out_rdata1,
  output [31:0] io_out_rdata2
);
  wire  regfile_clock; // @[regfile.scala 48:25]
  wire  regfile_reset; // @[regfile.scala 48:25]
  wire [4:0] regfile_rs1; // @[regfile.scala 48:25]
  wire [4:0] regfile_rs2; // @[regfile.scala 48:25]
  wire [4:0] regfile_rd; // @[regfile.scala 48:25]
  wire [31:0] regfile_wdata; // @[regfile.scala 48:25]
  wire  regfile_reg_wen; // @[regfile.scala 48:25]
  wire [31:0] regfile_rdata1; // @[regfile.scala 48:25]
  wire [31:0] regfile_rdata2; // @[regfile.scala 48:25]
  RegisterFileBB regfile ( // @[regfile.scala 48:25]
    .clock(regfile_clock),
    .reset(regfile_reset),
    .rs1(regfile_rs1),
    .rs2(regfile_rs2),
    .rd(regfile_rd),
    .wdata(regfile_wdata),
    .reg_wen(regfile_reg_wen),
    .rdata1(regfile_rdata1),
    .rdata2(regfile_rdata2)
  );
  assign io_out_rdata1 = regfile_rdata1; // @[regfile.scala 58:19]
  assign io_out_rdata2 = regfile_rdata2; // @[regfile.scala 59:19]
  assign regfile_clock = clock; // @[regfile.scala 50:24]
  assign regfile_reset = reset; // @[regfile.scala 51:24]
  assign regfile_rs1 = io_in_rs1; // @[regfile.scala 52:24]
  assign regfile_rs2 = io_in_rs2; // @[regfile.scala 53:24]
  assign regfile_rd = io_in_rd; // @[regfile.scala 54:24]
  assign regfile_wdata = io_in_wdata; // @[regfile.scala 55:24]
  assign regfile_reg_wen = io_in_reg_wen; // @[regfile.scala 56:24]
endmodule
module ISU(
  input         clock,
  input         reset,
  input         from_IDU_valid,
  input  [31:0] from_IDU_bits_imm,
  input  [31:0] from_IDU_bits_pc,
  input  [4:0]  from_IDU_bits_rs1,
  input  [4:0]  from_IDU_bits_rs2,
  input  [4:0]  from_IDU_bits_rd,
  input         from_IDU_bits_ctrl_sig_reg_wen,
  input  [2:0]  from_IDU_bits_ctrl_sig_fu_op,
  input         from_IDU_bits_ctrl_sig_mem_wen,
  input         from_IDU_bits_ctrl_sig_is_ebreak,
  input         from_IDU_bits_ctrl_sig_not_impl,
  input  [1:0]  from_IDU_bits_ctrl_sig_src1_op,
  input  [1:0]  from_IDU_bits_ctrl_sig_src2_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_alu_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_lsu_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_bru_op,
  input  [2:0]  from_IDU_bits_ctrl_sig_csr_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_mdu_op,
  input         from_WBU_bits_reg_wen,
  input  [31:0] from_WBU_bits_wdata,
  input  [4:0]  from_WBU_bits_rd,
  output        to_EXU_valid,
  output [31:0] to_EXU_bits_imm,
  output [31:0] to_EXU_bits_pc,
  output [31:0] to_EXU_bits_rdata1,
  output [31:0] to_EXU_bits_rdata2,
  output [4:0]  to_EXU_bits_rd,
  output        to_EXU_bits_ctrl_sig_reg_wen,
  output [2:0]  to_EXU_bits_ctrl_sig_fu_op,
  output        to_EXU_bits_ctrl_sig_mem_wen,
  output        to_EXU_bits_ctrl_sig_is_ebreak,
  output        to_EXU_bits_ctrl_sig_not_impl,
  output [1:0]  to_EXU_bits_ctrl_sig_src1_op,
  output [1:0]  to_EXU_bits_ctrl_sig_src2_op,
  output [3:0]  to_EXU_bits_ctrl_sig_alu_op,
  output [3:0]  to_EXU_bits_ctrl_sig_lsu_op,
  output [3:0]  to_EXU_bits_ctrl_sig_bru_op,
  output [2:0]  to_EXU_bits_ctrl_sig_csr_op,
  output [3:0]  to_EXU_bits_ctrl_sig_mdu_op
);
  wire  RegFile_i_clock; // @[ISU.scala 20:37]
  wire  RegFile_i_reset; // @[ISU.scala 20:37]
  wire [4:0] RegFile_i_io_in_rs1; // @[ISU.scala 20:37]
  wire [4:0] RegFile_i_io_in_rs2; // @[ISU.scala 20:37]
  wire [4:0] RegFile_i_io_in_rd; // @[ISU.scala 20:37]
  wire [31:0] RegFile_i_io_in_wdata; // @[ISU.scala 20:37]
  wire  RegFile_i_io_in_reg_wen; // @[ISU.scala 20:37]
  wire [31:0] RegFile_i_io_out_rdata1; // @[ISU.scala 20:37]
  wire [31:0] RegFile_i_io_out_rdata2; // @[ISU.scala 20:37]
  RegFile RegFile_i ( // @[ISU.scala 20:37]
    .clock(RegFile_i_clock),
    .reset(RegFile_i_reset),
    .io_in_rs1(RegFile_i_io_in_rs1),
    .io_in_rs2(RegFile_i_io_in_rs2),
    .io_in_rd(RegFile_i_io_in_rd),
    .io_in_wdata(RegFile_i_io_in_wdata),
    .io_in_reg_wen(RegFile_i_io_in_reg_wen),
    .io_out_rdata1(RegFile_i_io_out_rdata1),
    .io_out_rdata2(RegFile_i_io_out_rdata2)
  );
  assign to_EXU_valid = from_IDU_valid; // @[ISU.scala 18:20]
  assign to_EXU_bits_imm = from_IDU_bits_imm; // @[ISU.scala 33:26]
  assign to_EXU_bits_pc = from_IDU_bits_pc; // @[ISU.scala 34:26]
  assign to_EXU_bits_rdata1 = RegFile_i_io_out_rdata1; // @[ISU.scala 36:26]
  assign to_EXU_bits_rdata2 = RegFile_i_io_out_rdata2; // @[ISU.scala 37:26]
  assign to_EXU_bits_rd = from_IDU_bits_rd; // @[ISU.scala 35:26]
  assign to_EXU_bits_ctrl_sig_reg_wen = from_IDU_bits_ctrl_sig_reg_wen; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_fu_op = from_IDU_bits_ctrl_sig_fu_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_mem_wen = from_IDU_bits_ctrl_sig_mem_wen; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_is_ebreak = from_IDU_bits_ctrl_sig_is_ebreak; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_not_impl = from_IDU_bits_ctrl_sig_not_impl; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_src1_op = from_IDU_bits_ctrl_sig_src1_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_src2_op = from_IDU_bits_ctrl_sig_src2_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_alu_op = from_IDU_bits_ctrl_sig_alu_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_lsu_op = from_IDU_bits_ctrl_sig_lsu_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_bru_op = from_IDU_bits_ctrl_sig_bru_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_csr_op = from_IDU_bits_ctrl_sig_csr_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_mdu_op = from_IDU_bits_ctrl_sig_mdu_op; // @[ISU.scala 32:26]
  assign RegFile_i_clock = clock;
  assign RegFile_i_reset = reset;
  assign RegFile_i_io_in_rs1 = from_IDU_bits_rs1; // @[ISU.scala 24:29]
  assign RegFile_i_io_in_rs2 = from_IDU_bits_rs2; // @[ISU.scala 25:29]
  assign RegFile_i_io_in_rd = from_WBU_bits_rd; // @[ISU.scala 23:29]
  assign RegFile_i_io_in_wdata = from_WBU_bits_wdata; // @[ISU.scala 29:29]
  assign RegFile_i_io_in_reg_wen = from_WBU_bits_reg_wen; // @[ISU.scala 28:29]
endmodule
module Alu(
  input  [31:0] io_in_src1,
  input  [31:0] io_in_src2,
  input  [3:0]  io_in_op,
  output [31:0] io_out_result
);
  wire [4:0] shamt = io_in_src2[4:0]; // @[alu.scala 31:25]
  wire [31:0] _io_out_result_T_1 = io_in_src1 + io_in_src2; // @[alu.scala 36:42]
  wire [31:0] _io_out_result_T_3 = io_in_src1 - io_in_src2; // @[alu.scala 37:42]
  wire [31:0] _io_out_result_T_4 = io_in_src1 & io_in_src2; // @[alu.scala 38:42]
  wire [31:0] _io_out_result_T_5 = io_in_src1 | io_in_src2; // @[alu.scala 39:42]
  wire [31:0] _io_out_result_T_6 = io_in_src1 ^ io_in_src2; // @[alu.scala 40:42]
  wire  _io_out_result_T_9 = $signed(io_in_src1) < $signed(io_in_src2); // @[alu.scala 41:49]
  wire  _io_out_result_T_10 = io_in_src1 < io_in_src2; // @[alu.scala 42:42]
  wire [62:0] _GEN_0 = {{31'd0}, io_in_src1}; // @[alu.scala 43:42]
  wire [62:0] _io_out_result_T_11 = _GEN_0 << shamt; // @[alu.scala 43:42]
  wire [31:0] _io_out_result_T_12 = io_in_src1 >> shamt; // @[alu.scala 44:42]
  wire [31:0] _io_out_result_T_15 = $signed(io_in_src1) >>> shamt; // @[alu.scala 45:59]
  wire [31:0] _io_out_result_T_19 = 4'h1 == io_in_op ? _io_out_result_T_1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_21 = 4'h2 == io_in_op ? _io_out_result_T_3 : _io_out_result_T_19; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_23 = 4'h3 == io_in_op ? _io_out_result_T_4 : _io_out_result_T_21; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_25 = 4'h4 == io_in_op ? _io_out_result_T_5 : _io_out_result_T_23; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_27 = 4'h5 == io_in_op ? _io_out_result_T_6 : _io_out_result_T_25; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_29 = 4'h6 == io_in_op ? {{31'd0}, _io_out_result_T_9} : _io_out_result_T_27; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_31 = 4'h7 == io_in_op ? {{31'd0}, _io_out_result_T_10} : _io_out_result_T_29; // @[Mux.scala 81:58]
  wire [62:0] _io_out_result_T_33 = 4'h8 == io_in_op ? _io_out_result_T_11 : {{31'd0}, _io_out_result_T_31}; // @[Mux.scala 81:58]
  wire [62:0] _io_out_result_T_35 = 4'h9 == io_in_op ? {{31'd0}, _io_out_result_T_12} : _io_out_result_T_33; // @[Mux.scala 81:58]
  wire [62:0] _io_out_result_T_37 = 4'ha == io_in_op ? {{31'd0}, _io_out_result_T_15} : _io_out_result_T_35; // @[Mux.scala 81:58]
  assign io_out_result = _io_out_result_T_37[31:0]; // @[alu.scala 33:21]
endmodule
module Mdu(
  input  [31:0] io_in_src1,
  input  [31:0] io_in_src2,
  input  [3:0]  io_in_op,
  output [31:0] io_out_result
);
  wire [63:0] _io_out_result_T = io_in_src1 * io_in_src2; // @[mdu.scala 36:44]
  wire [63:0] _io_out_result_T_3 = $signed(io_in_src1) * $signed(io_in_src2); // @[mdu.scala 37:52]
  wire [31:0] _io_out_result_T_5 = _io_out_result_T_3[63:32]; // @[mdu.scala 37:86]
  wire [32:0] _io_out_result_T_7 = {1'b0,$signed(io_in_src2)}; // @[mdu.scala 38:52]
  wire [64:0] _io_out_result_T_8 = $signed(io_in_src1) * $signed(_io_out_result_T_7); // @[mdu.scala 38:52]
  wire [63:0] _io_out_result_T_10 = _io_out_result_T_8[63:0]; // @[mdu.scala 38:52]
  wire [31:0] _io_out_result_T_12 = _io_out_result_T_10[63:32]; // @[mdu.scala 38:79]
  wire [32:0] _io_out_result_T_18 = $signed(io_in_src1) / $signed(io_in_src2); // @[mdu.scala 40:70]
  wire [31:0] _io_out_result_T_19 = io_in_src1 / io_in_src2; // @[mdu.scala 41:44]
  wire [31:0] _io_out_result_T_23 = $signed(io_in_src1) % $signed(io_in_src2); // @[mdu.scala 42:70]
  wire [31:0] _io_out_result_T_24 = io_in_src1 % io_in_src2; // @[mdu.scala 43:44]
  wire [63:0] _io_out_result_T_28 = 4'h1 == io_in_op ? _io_out_result_T : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_30 = 4'h2 == io_in_op ? {{32'd0}, _io_out_result_T_5} : _io_out_result_T_28; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_32 = 4'h3 == io_in_op ? {{32'd0}, _io_out_result_T_12} : _io_out_result_T_30; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_34 = 4'h4 == io_in_op ? {{32'd0}, _io_out_result_T[63:32]} : _io_out_result_T_32; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_36 = 4'h5 == io_in_op ? {{31'd0}, _io_out_result_T_18} : _io_out_result_T_34; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_38 = 4'h6 == io_in_op ? {{32'd0}, _io_out_result_T_19} : _io_out_result_T_36; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_40 = 4'h7 == io_in_op ? {{32'd0}, _io_out_result_T_23} : _io_out_result_T_38; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_42 = 4'h8 == io_in_op ? {{32'd0}, _io_out_result_T_24} : _io_out_result_T_40; // @[Mux.scala 81:58]
  assign io_out_result = _io_out_result_T_42[31:0]; // @[mdu.scala 33:21]
endmodule
module Bru(
  input  [31:0] io_in_src1,
  input  [31:0] io_in_src2,
  input  [3:0]  io_in_op,
  output        io_out_ctrl_br
);
  wire  _io_out_ctrl_br_T = io_in_src1 == io_in_src2; // @[bru.scala 35:44]
  wire  _io_out_ctrl_br_T_1 = io_in_src1 != io_in_src2; // @[bru.scala 36:44]
  wire  _io_out_ctrl_br_T_4 = $signed(io_in_src1) < $signed(io_in_src2); // @[bru.scala 37:51]
  wire  _io_out_ctrl_br_T_7 = $signed(io_in_src1) >= $signed(io_in_src2); // @[bru.scala 38:51]
  wire  _io_out_ctrl_br_T_8 = io_in_src1 < io_in_src2; // @[bru.scala 39:51]
  wire  _io_out_ctrl_br_T_9 = io_in_src1 >= io_in_src2; // @[bru.scala 40:51]
  wire  _io_out_ctrl_br_T_15 = 4'h3 == io_in_op ? _io_out_ctrl_br_T : 4'h2 == io_in_op | 4'h1 == io_in_op; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_17 = 4'h4 == io_in_op ? _io_out_ctrl_br_T_1 : _io_out_ctrl_br_T_15; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_19 = 4'h5 == io_in_op ? _io_out_ctrl_br_T_4 : _io_out_ctrl_br_T_17; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_21 = 4'h6 == io_in_op ? _io_out_ctrl_br_T_7 : _io_out_ctrl_br_T_19; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_23 = 4'h7 == io_in_op ? _io_out_ctrl_br_T_8 : _io_out_ctrl_br_T_21; // @[Mux.scala 81:58]
  assign io_out_ctrl_br = 4'h8 == io_in_op ? _io_out_ctrl_br_T_9 : _io_out_ctrl_br_T_23; // @[Mux.scala 81:58]
endmodule
module Lsu(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_mem_wen,
  input  [31:0] io_in_addr,
  input  [31:0] io_in_wdata,
  input  [3:0]  io_in_op,
  output [31:0] io_out_rdata,
  output        io_out_end,
  output        io_out_idle,
  input         axi_ar_ready,
  output        axi_ar_valid,
  output [31:0] axi_ar_bits_addr,
  output        axi_r_ready,
  input         axi_r_valid,
  input  [31:0] axi_r_bits_data,
  input         axi_aw_ready,
  output        axi_aw_valid,
  output [31:0] axi_aw_bits_addr,
  input         axi_w_ready,
  output        axi_w_valid,
  output [31:0] axi_w_bits_data,
  output [3:0]  axi_w_bits_strb,
  output        axi_b_ready,
  input         axi_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[lsu.scala 35:24]
  wire  _state_T = axi_ar_ready & axi_ar_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_2 = axi_r_ready & axi_r_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_3 = _state_T_2 ? 3'h5 : 3'h2; // @[lsu.scala 53:25]
  wire  _state_T_4 = axi_aw_ready & axi_aw_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_5 = axi_w_ready & axi_w_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_7 = _state_T_4 & _state_T_5 ? 3'h4 : 3'h3; // @[lsu.scala 58:25]
  wire  _state_T_8 = axi_b_ready & axi_b_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_9 = _state_T_8 ? 3'h5 : 3'h4; // @[lsu.scala 61:25]
  wire [2:0] _GEN_2 = 3'h5 == state ? 3'h0 : state; // @[lsu.scala 36:20 64:19 35:24]
  wire [2:0] _GEN_3 = 3'h4 == state ? _state_T_9 : _GEN_2; // @[lsu.scala 36:20 61:19]
  wire [2:0] _GEN_4 = 3'h3 == state ? _state_T_7 : _GEN_3; // @[lsu.scala 36:20 58:19]
  wire [1:0] addr_low_2 = io_in_addr[1:0]; // @[lsu.scala 71:31]
  wire [23:0] _lb_rdata_T_2 = axi_r_bits_data[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_4 = {_lb_rdata_T_2,axi_r_bits_data[7:0]}; // @[Cat.scala 33:92]
  wire [23:0] _lb_rdata_T_7 = axi_r_bits_data[15] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_9 = {_lb_rdata_T_7,axi_r_bits_data[15:8]}; // @[Cat.scala 33:92]
  wire [23:0] _lb_rdata_T_12 = axi_r_bits_data[23] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_14 = {_lb_rdata_T_12,axi_r_bits_data[23:16]}; // @[Cat.scala 33:92]
  wire [23:0] _lb_rdata_T_17 = axi_r_bits_data[31] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_19 = {_lb_rdata_T_17,axi_r_bits_data[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _lb_rdata_T_21 = 2'h1 == addr_low_2 ? _lb_rdata_T_9 : _lb_rdata_T_4; // @[Mux.scala 81:58]
  wire [31:0] _lb_rdata_T_23 = 2'h2 == addr_low_2 ? _lb_rdata_T_14 : _lb_rdata_T_21; // @[Mux.scala 81:58]
  wire [31:0] lb_rdata = 2'h3 == addr_low_2 ? _lb_rdata_T_19 : _lb_rdata_T_23; // @[Mux.scala 81:58]
  wire [31:0] _lbu_rdata_T_2 = {24'h0,axi_r_bits_data[7:0]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_5 = {24'h0,axi_r_bits_data[15:8]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_8 = {24'h0,axi_r_bits_data[23:16]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_11 = {24'h0,axi_r_bits_data[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_13 = 2'h1 == addr_low_2 ? _lbu_rdata_T_5 : _lbu_rdata_T_2; // @[Mux.scala 81:58]
  wire [31:0] _lbu_rdata_T_15 = 2'h2 == addr_low_2 ? _lbu_rdata_T_8 : _lbu_rdata_T_13; // @[Mux.scala 81:58]
  wire [31:0] lbu_rdata = 2'h3 == addr_low_2 ? _lbu_rdata_T_11 : _lbu_rdata_T_15; // @[Mux.scala 81:58]
  wire [15:0] _lh_rdata_T_2 = axi_r_bits_data[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lh_rdata_T_4 = {_lh_rdata_T_2,axi_r_bits_data[15:0]}; // @[Cat.scala 33:92]
  wire [15:0] _lh_rdata_T_7 = axi_r_bits_data[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lh_rdata_T_9 = {_lh_rdata_T_7,axi_r_bits_data[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _lh_rdata_T_11 = 2'h0 == addr_low_2 ? _lh_rdata_T_4 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] lh_rdata = 2'h2 == addr_low_2 ? _lh_rdata_T_9 : _lh_rdata_T_11; // @[Mux.scala 81:58]
  wire [31:0] _lhu_rdata_T_2 = {16'h0,axi_r_bits_data[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _lhu_rdata_T_5 = {16'h0,axi_r_bits_data[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _lhu_rdata_T_7 = 2'h0 == addr_low_2 ? _lhu_rdata_T_2 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] lhu_rdata = 2'h2 == addr_low_2 ? _lhu_rdata_T_5 : _lhu_rdata_T_7; // @[Mux.scala 81:58]
  wire [1:0] _sb_wmask_T_1 = 2'h1 == addr_low_2 ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [2:0] _sb_wmask_T_3 = 2'h2 == addr_low_2 ? 3'h4 : {{1'd0}, _sb_wmask_T_1}; // @[Mux.scala 81:58]
  wire [3:0] sb_wmask = 2'h3 == addr_low_2 ? 4'h8 : {{1'd0}, _sb_wmask_T_3}; // @[Mux.scala 81:58]
  wire [1:0] _sh_wmask_T_1 = 2'h0 == addr_low_2 ? 2'h3 : 2'h0; // @[Mux.scala 81:58]
  wire [3:0] sh_wmask = 2'h2 == addr_low_2 ? 4'hc : {{2'd0}, _sh_wmask_T_1}; // @[Mux.scala 81:58]
  wire [3:0] _wmask_T_1 = 4'h6 == io_in_op ? sb_wmask : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _wmask_T_3 = 4'h7 == io_in_op ? sh_wmask : _wmask_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_3 = 4'h1 == io_in_op ? lb_rdata : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_5 = 4'h4 == io_in_op ? lbu_rdata : _io_out_rdata_T_3; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_7 = 4'h2 == io_in_op ? lh_rdata : _io_out_rdata_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_9 = 4'h5 == io_in_op ? lhu_rdata : _io_out_rdata_T_7; // @[Mux.scala 81:58]
  assign io_out_rdata = 4'h3 == io_in_op ? axi_r_bits_data : _io_out_rdata_T_9; // @[Mux.scala 81:58]
  assign io_out_end = 3'h5 == state; // @[Mux.scala 81:61]
  assign io_out_idle = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_ar_valid = 3'h1 == state; // @[Mux.scala 81:61]
  assign axi_ar_bits_addr = io_in_addr; // @[lsu.scala 148:22]
  assign axi_r_ready = 3'h2 == state; // @[Mux.scala 81:61]
  assign axi_aw_valid = 3'h3 == state; // @[Mux.scala 81:61]
  assign axi_aw_bits_addr = io_in_addr; // @[lsu.scala 151:22]
  assign axi_w_valid = 3'h3 == state; // @[Mux.scala 81:61]
  assign axi_w_bits_data = io_in_wdata; // @[lsu.scala 153:22]
  assign axi_w_bits_strb = 4'h8 == io_in_op ? 4'hf : _wmask_T_3; // @[Mux.scala 81:58]
  assign axi_b_ready = 3'h4 == state; // @[Mux.scala 81:61]
  always @(posedge clock) begin
    if (reset) begin // @[lsu.scala 35:24]
      state <= 3'h0; // @[lsu.scala 35:24]
    end else if (3'h0 == state) begin // @[lsu.scala 36:20]
      if (io_in_valid) begin // @[lsu.scala 38:32]
        if (io_in_mem_wen) begin // @[lsu.scala 39:38]
          state <= 3'h3; // @[lsu.scala 40:27]
        end else begin
          state <= 3'h1; // @[lsu.scala 42:27]
        end
      end else begin
        state <= 3'h0; // @[lsu.scala 45:23]
      end
    end else if (3'h1 == state) begin // @[lsu.scala 36:20]
      if (_state_T) begin // @[lsu.scala 50:25]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[lsu.scala 36:20]
      state <= _state_T_3; // @[lsu.scala 53:19]
    end else begin
      state <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csr(
  input         clock,
  input         reset,
  input  [2:0]  io_in_op,
  input  [31:0] io_in_cur_pc,
  input  [31:0] io_in_csr_id,
  input  [31:0] io_in_wdata,
  output        io_out_csr_br,
  output [31:0] io_out_csr_addr,
  output [31:0] io_out_r_csr,
  output [31:0] io_out_difftest_mcause,
  output [31:0] io_out_difftest_mepc,
  output [31:0] io_out_difftest_mstatus,
  output [31:0] io_out_difftest_mtvec
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_mepc; // @[csr.scala 32:28]
  reg [31:0] reg_mcause; // @[csr.scala 33:28]
  reg [31:0] reg_mstatus; // @[csr.scala 34:28]
  reg [31:0] reg_mtvec; // @[csr.scala 35:28]
  wire [31:0] _reg_mcause_csrrs_T = io_in_wdata | reg_mcause; // @[csr.scala 51:32]
  wire [31:0] _reg_mepc_csrrs_T = io_in_wdata | reg_mepc; // @[csr.scala 63:30]
  wire [31:0] _reg_mstatus_csrrs_T = io_in_wdata | reg_mstatus; // @[csr.scala 75:33]
  wire [31:0] _reg_mstatus_T_5 = {reg_mstatus[31:13],2'h3,reg_mstatus[10:8],reg_mstatus[3],reg_mstatus[6:4],1'h0,
    reg_mstatus[2:0]}; // @[Cat.scala 33:92]
  wire [30:0] _reg_mstatus_T_11 = {reg_mstatus[31:13],1'h0,reg_mstatus[10:8],1'h1,reg_mstatus[6:4],reg_mstatus[7],
    reg_mstatus[2:0]}; // @[Cat.scala 33:92]
  wire [31:0] _reg_mstatus_T_13 = 3'h1 == io_in_op ? _reg_mstatus_T_5 : reg_mstatus; // @[Mux.scala 81:58]
  wire [31:0] _reg_mtvec_csrrs_T = io_in_wdata | reg_mtvec; // @[csr.scala 100:31]
  wire [31:0] _io_out_csr_addr_T_1 = 3'h1 == io_in_op ? reg_mtvec : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_r_csr_T_1 = 32'h305 == io_in_csr_id ? reg_mtvec : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_r_csr_T_3 = 32'h341 == io_in_csr_id ? reg_mepc : _io_out_r_csr_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_out_r_csr_T_5 = 32'h342 == io_in_csr_id ? reg_mcause : _io_out_r_csr_T_3; // @[Mux.scala 81:58]
  assign io_out_csr_br = 3'h2 == io_in_op | 3'h1 == io_in_op; // @[Mux.scala 81:58]
  assign io_out_csr_addr = 3'h2 == io_in_op ? reg_mepc : _io_out_csr_addr_T_1; // @[Mux.scala 81:58]
  assign io_out_r_csr = 32'h300 == io_in_csr_id ? reg_mstatus : _io_out_r_csr_T_5; // @[Mux.scala 81:58]
  assign io_out_difftest_mcause = reg_mcause; // @[csr.scala 125:27]
  assign io_out_difftest_mepc = reg_mepc; // @[csr.scala 126:27]
  assign io_out_difftest_mstatus = reg_mstatus; // @[csr.scala 127:27]
  assign io_out_difftest_mtvec = reg_mtvec; // @[csr.scala 128:27]
  always @(posedge clock) begin
    if (reset) begin // @[csr.scala 32:28]
      reg_mepc <= 32'h0; // @[csr.scala 32:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h341 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mepc <= _reg_mepc_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h341 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mepc <= io_in_wdata;
      end
    end else if (3'h1 == io_in_op) begin // @[Mux.scala 81:58]
      reg_mepc <= io_in_cur_pc;
    end
    if (reset) begin // @[csr.scala 33:28]
      reg_mcause <= 32'h0; // @[csr.scala 33:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h342 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mcause <= _reg_mcause_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h342 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mcause <= io_in_wdata;
      end
    end else if (3'h1 == io_in_op) begin // @[Mux.scala 81:58]
      reg_mcause <= 32'hb;
    end
    if (reset) begin // @[csr.scala 34:28]
      reg_mstatus <= 32'h0; // @[csr.scala 34:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h300 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mstatus <= _reg_mstatus_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h300 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mstatus <= io_in_wdata;
      end
    end else if (3'h2 == io_in_op) begin // @[Mux.scala 81:58]
      reg_mstatus <= {{1'd0}, _reg_mstatus_T_11};
    end else begin
      reg_mstatus <= _reg_mstatus_T_13;
    end
    if (reset) begin // @[csr.scala 35:28]
      reg_mtvec <= 32'h0; // @[csr.scala 35:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h305 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mtvec <= _reg_mtvec_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h305 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mtvec <= io_in_wdata;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mepc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mcause = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_mtvec = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ebreak_moudle(
  input   is_ebreak
);
  wire  EbreakBB_i1_is_ebreak; // @[ebreak.scala 21:29]
  EbreakBB EbreakBB_i1 ( // @[ebreak.scala 21:29]
    .is_ebreak(EbreakBB_i1_is_ebreak)
  );
  assign EbreakBB_i1_is_ebreak = is_ebreak; // @[ebreak.scala 23:30]
endmodule
module not_impl_moudle(
  input   not_impl
);
  wire  NotImplBB_i1_not_impl; // @[not_impl.scala 21:30]
  NotImplBB NotImplBB_i1 ( // @[not_impl.scala 21:30]
    .not_impl(NotImplBB_i1_not_impl)
  );
  assign NotImplBB_i1_not_impl = not_impl; // @[not_impl.scala 23:30]
endmodule
module EXU(
  input         clock,
  input         reset,
  output        from_ISU_ready,
  input         from_ISU_valid,
  input  [31:0] from_ISU_bits_imm,
  input  [31:0] from_ISU_bits_pc,
  input  [31:0] from_ISU_bits_rdata1,
  input  [31:0] from_ISU_bits_rdata2,
  input  [4:0]  from_ISU_bits_rd,
  input         from_ISU_bits_ctrl_sig_reg_wen,
  input  [2:0]  from_ISU_bits_ctrl_sig_fu_op,
  input         from_ISU_bits_ctrl_sig_mem_wen,
  input         from_ISU_bits_ctrl_sig_is_ebreak,
  input         from_ISU_bits_ctrl_sig_not_impl,
  input  [1:0]  from_ISU_bits_ctrl_sig_src1_op,
  input  [1:0]  from_ISU_bits_ctrl_sig_src2_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_alu_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_lsu_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_bru_op,
  input  [2:0]  from_ISU_bits_ctrl_sig_csr_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_mdu_op,
  output        to_WBU_valid,
  output [31:0] to_WBU_bits_alu_result,
  output [31:0] to_WBU_bits_mdu_result,
  output [31:0] to_WBU_bits_lsu_rdata,
  output [31:0] to_WBU_bits_csr_rdata,
  output [31:0] to_WBU_bits_pc,
  output        to_WBU_bits_reg_wen,
  output [4:0]  to_WBU_bits_rd,
  output [2:0]  to_WBU_bits_fu_op,
  output        to_IFU_bits_bru_ctrl_br,
  output [31:0] to_IFU_bits_bru_addr,
  output        to_IFU_bits_csr_ctrl_br,
  output [31:0] to_IFU_bits_csr_addr,
  output [31:0] difftest_mcause,
  output [31:0] difftest_mepc,
  output [31:0] difftest_mstatus,
  output [31:0] difftest_mtvec,
  input         lsu_axi_master_ar_ready,
  output        lsu_axi_master_ar_valid,
  output [31:0] lsu_axi_master_ar_bits_addr,
  output        lsu_axi_master_r_ready,
  input         lsu_axi_master_r_valid,
  input  [31:0] lsu_axi_master_r_bits_data,
  input         lsu_axi_master_aw_ready,
  output        lsu_axi_master_aw_valid,
  output [31:0] lsu_axi_master_aw_bits_addr,
  input         lsu_axi_master_w_ready,
  output        lsu_axi_master_w_valid,
  output [31:0] lsu_axi_master_w_bits_data,
  output [3:0]  lsu_axi_master_w_bits_strb,
  output        lsu_axi_master_b_ready,
  input         lsu_axi_master_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] Alu_i_io_in_src1; // @[EXU.scala 22:37]
  wire [31:0] Alu_i_io_in_src2; // @[EXU.scala 22:37]
  wire [3:0] Alu_i_io_in_op; // @[EXU.scala 22:37]
  wire [31:0] Alu_i_io_out_result; // @[EXU.scala 22:37]
  wire [31:0] Mdu_i_io_in_src1; // @[EXU.scala 23:37]
  wire [31:0] Mdu_i_io_in_src2; // @[EXU.scala 23:37]
  wire [3:0] Mdu_i_io_in_op; // @[EXU.scala 23:37]
  wire [31:0] Mdu_i_io_out_result; // @[EXU.scala 23:37]
  wire [31:0] Bru_i_io_in_src1; // @[EXU.scala 24:37]
  wire [31:0] Bru_i_io_in_src2; // @[EXU.scala 24:37]
  wire [3:0] Bru_i_io_in_op; // @[EXU.scala 24:37]
  wire  Bru_i_io_out_ctrl_br; // @[EXU.scala 24:37]
  wire  Lsu_i_clock; // @[EXU.scala 25:37]
  wire  Lsu_i_reset; // @[EXU.scala 25:37]
  wire  Lsu_i_io_in_valid; // @[EXU.scala 25:37]
  wire  Lsu_i_io_in_mem_wen; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_io_in_addr; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_io_in_wdata; // @[EXU.scala 25:37]
  wire [3:0] Lsu_i_io_in_op; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_io_out_rdata; // @[EXU.scala 25:37]
  wire  Lsu_i_io_out_end; // @[EXU.scala 25:37]
  wire  Lsu_i_io_out_idle; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_ar_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_ar_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_ar_bits_addr; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_r_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_r_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_r_bits_data; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_aw_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_aw_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_aw_bits_addr; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_w_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_w_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_w_bits_data; // @[EXU.scala 25:37]
  wire [3:0] Lsu_i_axi_w_bits_strb; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_b_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_b_valid; // @[EXU.scala 25:37]
  wire  Csr_i_clock; // @[EXU.scala 26:37]
  wire  Csr_i_reset; // @[EXU.scala 26:37]
  wire [2:0] Csr_i_io_in_op; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_in_cur_pc; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_in_csr_id; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_in_wdata; // @[EXU.scala 26:37]
  wire  Csr_i_io_out_csr_br; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_csr_addr; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_r_csr; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mcause; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mepc; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mstatus; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mtvec; // @[EXU.scala 26:37]
  wire  ebreak_moudle_i_is_ebreak; // @[EXU.scala 27:37]
  wire  not_impl_moudle_i_not_impl; // @[EXU.scala 28:37]
  reg [1:0] state; // @[EXU.scala 37:24]
  wire  _state_T = from_ISU_ready & from_ISU_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_T_2 = Lsu_i_io_out_idle ? 2'h2 : 2'h1; // @[EXU.scala 45:29]
  wire [1:0] _state_T_3 = Lsu_i_io_out_end ? 2'h3 : 2'h2; // @[EXU.scala 51:25]
  wire [1:0] _GEN_1 = 2'h3 == state ? 2'h0 : state; // @[EXU.scala 38:20 54:19 37:24]
  wire [31:0] _Alu_i_io_in_src1_T_1 = 2'h2 == from_ISU_bits_ctrl_sig_src1_op ? from_ISU_bits_rdata1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _Alu_i_io_in_src2_T_1 = 2'h2 == from_ISU_bits_ctrl_sig_src2_op ? from_ISU_bits_rdata2 : 32'h0; // @[Mux.scala 81:58]
  Alu Alu_i ( // @[EXU.scala 22:37]
    .io_in_src1(Alu_i_io_in_src1),
    .io_in_src2(Alu_i_io_in_src2),
    .io_in_op(Alu_i_io_in_op),
    .io_out_result(Alu_i_io_out_result)
  );
  Mdu Mdu_i ( // @[EXU.scala 23:37]
    .io_in_src1(Mdu_i_io_in_src1),
    .io_in_src2(Mdu_i_io_in_src2),
    .io_in_op(Mdu_i_io_in_op),
    .io_out_result(Mdu_i_io_out_result)
  );
  Bru Bru_i ( // @[EXU.scala 24:37]
    .io_in_src1(Bru_i_io_in_src1),
    .io_in_src2(Bru_i_io_in_src2),
    .io_in_op(Bru_i_io_in_op),
    .io_out_ctrl_br(Bru_i_io_out_ctrl_br)
  );
  Lsu Lsu_i ( // @[EXU.scala 25:37]
    .clock(Lsu_i_clock),
    .reset(Lsu_i_reset),
    .io_in_valid(Lsu_i_io_in_valid),
    .io_in_mem_wen(Lsu_i_io_in_mem_wen),
    .io_in_addr(Lsu_i_io_in_addr),
    .io_in_wdata(Lsu_i_io_in_wdata),
    .io_in_op(Lsu_i_io_in_op),
    .io_out_rdata(Lsu_i_io_out_rdata),
    .io_out_end(Lsu_i_io_out_end),
    .io_out_idle(Lsu_i_io_out_idle),
    .axi_ar_ready(Lsu_i_axi_ar_ready),
    .axi_ar_valid(Lsu_i_axi_ar_valid),
    .axi_ar_bits_addr(Lsu_i_axi_ar_bits_addr),
    .axi_r_ready(Lsu_i_axi_r_ready),
    .axi_r_valid(Lsu_i_axi_r_valid),
    .axi_r_bits_data(Lsu_i_axi_r_bits_data),
    .axi_aw_ready(Lsu_i_axi_aw_ready),
    .axi_aw_valid(Lsu_i_axi_aw_valid),
    .axi_aw_bits_addr(Lsu_i_axi_aw_bits_addr),
    .axi_w_ready(Lsu_i_axi_w_ready),
    .axi_w_valid(Lsu_i_axi_w_valid),
    .axi_w_bits_data(Lsu_i_axi_w_bits_data),
    .axi_w_bits_strb(Lsu_i_axi_w_bits_strb),
    .axi_b_ready(Lsu_i_axi_b_ready),
    .axi_b_valid(Lsu_i_axi_b_valid)
  );
  Csr Csr_i ( // @[EXU.scala 26:37]
    .clock(Csr_i_clock),
    .reset(Csr_i_reset),
    .io_in_op(Csr_i_io_in_op),
    .io_in_cur_pc(Csr_i_io_in_cur_pc),
    .io_in_csr_id(Csr_i_io_in_csr_id),
    .io_in_wdata(Csr_i_io_in_wdata),
    .io_out_csr_br(Csr_i_io_out_csr_br),
    .io_out_csr_addr(Csr_i_io_out_csr_addr),
    .io_out_r_csr(Csr_i_io_out_r_csr),
    .io_out_difftest_mcause(Csr_i_io_out_difftest_mcause),
    .io_out_difftest_mepc(Csr_i_io_out_difftest_mepc),
    .io_out_difftest_mstatus(Csr_i_io_out_difftest_mstatus),
    .io_out_difftest_mtvec(Csr_i_io_out_difftest_mtvec)
  );
  ebreak_moudle ebreak_moudle_i ( // @[EXU.scala 27:37]
    .is_ebreak(ebreak_moudle_i_is_ebreak)
  );
  not_impl_moudle not_impl_moudle_i ( // @[EXU.scala 28:37]
    .not_impl(not_impl_moudle_i_not_impl)
  );
  assign from_ISU_ready = 2'h0 == state; // @[Mux.scala 81:61]
  assign to_WBU_valid = 2'h3 == state; // @[Mux.scala 81:61]
  assign to_WBU_bits_alu_result = Alu_i_io_out_result; // @[EXU.scala 102:28]
  assign to_WBU_bits_mdu_result = Mdu_i_io_out_result; // @[EXU.scala 103:28]
  assign to_WBU_bits_lsu_rdata = Lsu_i_io_out_rdata; // @[EXU.scala 104:28]
  assign to_WBU_bits_csr_rdata = Csr_i_io_out_r_csr; // @[EXU.scala 105:28]
  assign to_WBU_bits_pc = from_ISU_bits_pc; // @[EXU.scala 107:28]
  assign to_WBU_bits_reg_wen = from_ISU_bits_ctrl_sig_reg_wen; // @[EXU.scala 108:28]
  assign to_WBU_bits_rd = from_ISU_bits_rd; // @[EXU.scala 110:28]
  assign to_WBU_bits_fu_op = from_ISU_bits_ctrl_sig_fu_op; // @[EXU.scala 109:28]
  assign to_IFU_bits_bru_ctrl_br = Bru_i_io_out_ctrl_br; // @[EXU.scala 112:33]
  assign to_IFU_bits_bru_addr = Alu_i_io_out_result; // @[EXU.scala 113:33]
  assign to_IFU_bits_csr_ctrl_br = Csr_i_io_out_csr_br; // @[EXU.scala 114:33]
  assign to_IFU_bits_csr_addr = Csr_i_io_out_csr_addr; // @[EXU.scala 115:33]
  assign difftest_mcause = Csr_i_io_out_difftest_mcause; // @[EXU.scala 117:14]
  assign difftest_mepc = Csr_i_io_out_difftest_mepc; // @[EXU.scala 117:14]
  assign difftest_mstatus = Csr_i_io_out_difftest_mstatus; // @[EXU.scala 117:14]
  assign difftest_mtvec = Csr_i_io_out_difftest_mtvec; // @[EXU.scala 117:14]
  assign lsu_axi_master_ar_valid = Lsu_i_axi_ar_valid; // @[EXU.scala 118:20]
  assign lsu_axi_master_ar_bits_addr = Lsu_i_axi_ar_bits_addr; // @[EXU.scala 118:20]
  assign lsu_axi_master_r_ready = Lsu_i_axi_r_ready; // @[EXU.scala 118:20]
  assign lsu_axi_master_aw_valid = Lsu_i_axi_aw_valid; // @[EXU.scala 118:20]
  assign lsu_axi_master_aw_bits_addr = Lsu_i_axi_aw_bits_addr; // @[EXU.scala 118:20]
  assign lsu_axi_master_w_valid = Lsu_i_axi_w_valid; // @[EXU.scala 118:20]
  assign lsu_axi_master_w_bits_data = Lsu_i_axi_w_bits_data; // @[EXU.scala 118:20]
  assign lsu_axi_master_w_bits_strb = Lsu_i_axi_w_bits_strb; // @[EXU.scala 118:20]
  assign lsu_axi_master_b_ready = Lsu_i_axi_b_ready; // @[EXU.scala 118:20]
  assign Alu_i_io_in_src1 = 2'h1 == from_ISU_bits_ctrl_sig_src1_op ? from_ISU_bits_pc : _Alu_i_io_in_src1_T_1; // @[Mux.scala 81:58]
  assign Alu_i_io_in_src2 = 2'h3 == from_ISU_bits_ctrl_sig_src2_op ? from_ISU_bits_imm : _Alu_i_io_in_src2_T_1; // @[Mux.scala 81:58]
  assign Alu_i_io_in_op = from_ISU_bits_ctrl_sig_alu_op; // @[EXU.scala 62:20]
  assign Mdu_i_io_in_src1 = from_ISU_bits_rdata1; // @[EXU.scala 74:24]
  assign Mdu_i_io_in_src2 = from_ISU_bits_rdata2; // @[EXU.scala 75:24]
  assign Mdu_i_io_in_op = from_ISU_bits_ctrl_sig_mdu_op; // @[EXU.scala 73:24]
  assign Bru_i_io_in_src1 = from_ISU_bits_rdata1; // @[EXU.scala 87:24]
  assign Bru_i_io_in_src2 = from_ISU_bits_rdata2; // @[EXU.scala 88:24]
  assign Bru_i_io_in_op = from_ISU_bits_ctrl_sig_bru_op; // @[EXU.scala 86:24]
  assign Lsu_i_clock = clock;
  assign Lsu_i_reset = reset;
  assign Lsu_i_io_in_valid = 2'h2 == state; // @[Mux.scala 81:61]
  assign Lsu_i_io_in_mem_wen = from_ISU_bits_ctrl_sig_mem_wen; // @[EXU.scala 80:25]
  assign Lsu_i_io_in_addr = Alu_i_io_out_result; // @[EXU.scala 78:25]
  assign Lsu_i_io_in_wdata = from_ISU_bits_rdata2; // @[EXU.scala 79:25]
  assign Lsu_i_io_in_op = from_ISU_bits_ctrl_sig_lsu_op; // @[EXU.scala 81:25]
  assign Lsu_i_axi_ar_ready = lsu_axi_master_ar_ready; // @[EXU.scala 118:20]
  assign Lsu_i_axi_r_valid = lsu_axi_master_r_valid; // @[EXU.scala 118:20]
  assign Lsu_i_axi_r_bits_data = lsu_axi_master_r_bits_data; // @[EXU.scala 118:20]
  assign Lsu_i_axi_aw_ready = lsu_axi_master_aw_ready; // @[EXU.scala 118:20]
  assign Lsu_i_axi_w_ready = lsu_axi_master_w_ready; // @[EXU.scala 118:20]
  assign Lsu_i_axi_b_valid = lsu_axi_master_b_valid; // @[EXU.scala 118:20]
  assign Csr_i_clock = clock;
  assign Csr_i_reset = reset;
  assign Csr_i_io_in_op = from_ISU_bits_ctrl_sig_csr_op; // @[EXU.scala 91:25]
  assign Csr_i_io_in_cur_pc = from_ISU_bits_pc; // @[EXU.scala 92:25]
  assign Csr_i_io_in_csr_id = from_ISU_bits_imm; // @[EXU.scala 93:25]
  assign Csr_i_io_in_wdata = from_ISU_bits_rdata1; // @[EXU.scala 95:25]
  assign ebreak_moudle_i_is_ebreak = from_ISU_bits_ctrl_sig_is_ebreak; // @[EXU.scala 98:32]
  assign not_impl_moudle_i_not_impl = from_ISU_bits_ctrl_sig_not_impl; // @[EXU.scala 100:32]
  always @(posedge clock) begin
    if (reset) begin // @[EXU.scala 37:24]
      state <= 2'h0; // @[EXU.scala 37:24]
    end else if (2'h0 == state) begin // @[EXU.scala 38:20]
      if (_state_T) begin // @[EXU.scala 40:25]
        state <= 2'h1;
      end else begin
        state <= 2'h0;
      end
    end else if (2'h1 == state) begin // @[EXU.scala 38:20]
      if (from_ISU_bits_ctrl_sig_fu_op == 3'h4) begin // @[EXU.scala 44:69]
        state <= _state_T_2; // @[EXU.scala 45:23]
      end else begin
        state <= 2'h3; // @[EXU.scala 47:23]
      end
    end else if (2'h2 == state) begin // @[EXU.scala 38:20]
      state <= _state_T_3; // @[EXU.scala 51:19]
    end else begin
      state <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  output        from_EXU_ready,
  input         from_EXU_valid,
  input  [31:0] from_EXU_bits_alu_result,
  input  [31:0] from_EXU_bits_mdu_result,
  input  [31:0] from_EXU_bits_lsu_rdata,
  input  [31:0] from_EXU_bits_csr_rdata,
  input  [31:0] from_EXU_bits_pc,
  input         from_EXU_bits_reg_wen,
  input  [4:0]  from_EXU_bits_rd,
  input  [2:0]  from_EXU_bits_fu_op,
  output        to_ISU_bits_reg_wen,
  output [31:0] to_ISU_bits_wdata,
  output [4:0]  to_ISU_bits_rd,
  output        to_IFU_valid
);
  wire  _to_ISU_bits_reg_wen_T = from_EXU_ready & from_EXU_valid; // @[Decoupled.scala 51:35]
  wire [31:0] _to_ISU_bits_wdata_T_1 = from_EXU_bits_pc + 32'h4; // @[WBU.scala 25:47]
  wire [31:0] _to_ISU_bits_wdata_T_3 = 3'h1 == from_EXU_bits_fu_op ? from_EXU_bits_alu_result : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_wdata_T_5 = 3'h4 == from_EXU_bits_fu_op ? from_EXU_bits_lsu_rdata : _to_ISU_bits_wdata_T_3; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_wdata_T_7 = 3'h3 == from_EXU_bits_fu_op ? _to_ISU_bits_wdata_T_1 : _to_ISU_bits_wdata_T_5; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_wdata_T_9 = 3'h5 == from_EXU_bits_fu_op ? from_EXU_bits_csr_rdata : _to_ISU_bits_wdata_T_7; // @[Mux.scala 81:58]
  assign from_EXU_ready = 1'h1; // @[WBU.scala 14:20]
  assign to_ISU_bits_reg_wen = _to_ISU_bits_reg_wen_T & from_EXU_bits_reg_wen; // @[WBU.scala 19:31]
  assign to_ISU_bits_wdata = 3'h2 == from_EXU_bits_fu_op ? from_EXU_bits_mdu_result : _to_ISU_bits_wdata_T_9; // @[Mux.scala 81:58]
  assign to_ISU_bits_rd = from_EXU_bits_rd; // @[WBU.scala 20:25]
  assign to_IFU_valid = from_EXU_valid; // @[WBU.scala 16:20]
endmodule
module IFU_cache(
  input         clock,
  input         reset,
  output        to_IDU_valid,
  output [31:0] to_IDU_bits_inst,
  output [31:0] to_IDU_bits_pc,
  input         from_EXU_bits_bru_ctrl_br,
  input  [31:0] from_EXU_bits_bru_addr,
  input         from_EXU_bits_csr_ctrl_br,
  input  [31:0] from_EXU_bits_csr_addr,
  output        from_WBU_ready,
  input         from_WBU_valid,
  input         to_cache_ready,
  output        to_cache_valid,
  output [31:0] to_cache_bits_addr,
  output        from_cache_ready,
  input         from_cache_valid,
  input  [31:0] from_cache_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_PC; // @[IFU.scala 148:26]
  wire [31:0] _next_PC_T_1 = reg_PC + 32'h4; // @[IFU.scala 156:27]
  wire  _reg_PC_T = from_WBU_ready & from_WBU_valid; // @[Decoupled.scala 51:35]
  reg [1:0] state_ifu; // @[IFU.scala 164:28]
  wire  _state_ifu_T = to_cache_ready & to_cache_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_ifu_T_1 = _state_ifu_T ? 2'h1 : 2'h0; // @[IFU.scala 166:26]
  wire  _state_ifu_T_2 = from_cache_ready & from_cache_valid; // @[Decoupled.scala 51:35]
  assign to_IDU_valid = 2'h2 == state_ifu; // @[Mux.scala 81:61]
  assign to_IDU_bits_inst = to_IDU_valid ? from_cache_bits_data : 32'h13; // @[IFU.scala 178:28]
  assign to_IDU_bits_pc = reg_PC; // @[IFU.scala 179:22]
  assign from_WBU_ready = 2'h2 == state_ifu; // @[Mux.scala 81:61]
  assign to_cache_valid = 2'h0 == state_ifu; // @[Mux.scala 81:61]
  assign to_cache_bits_addr = reg_PC; // @[IFU.scala 173:24]
  assign from_cache_ready = 2'h1 == state_ifu; // @[Mux.scala 81:61]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 148:26]
      reg_PC <= 32'h80000000; // @[IFU.scala 148:26]
    end else if (_reg_PC_T) begin // @[IFU.scala 160:18]
      if (from_EXU_bits_bru_ctrl_br) begin // @[IFU.scala 151:38]
        reg_PC <= from_EXU_bits_bru_addr; // @[IFU.scala 152:17]
      end else if (from_EXU_bits_csr_ctrl_br) begin // @[IFU.scala 153:45]
        reg_PC <= from_EXU_bits_csr_addr; // @[IFU.scala 154:17]
      end else begin
        reg_PC <= _next_PC_T_1; // @[IFU.scala 156:17]
      end
    end
    if (reset) begin // @[IFU.scala 164:28]
      state_ifu <= 2'h0; // @[IFU.scala 164:28]
    end else if (2'h2 == state_ifu) begin // @[Mux.scala 81:58]
      if (_reg_PC_T) begin // @[IFU.scala 168:28]
        state_ifu <= 2'h0;
      end else begin
        state_ifu <= 2'h2;
      end
    end else if (2'h1 == state_ifu) begin // @[Mux.scala 81:58]
      if (_state_ifu_T_2) begin // @[IFU.scala 167:28]
        state_ifu <= 2'h2;
      end else begin
        state_ifu <= 2'h1;
      end
    end else if (2'h0 == state_ifu) begin // @[Mux.scala 81:58]
      state_ifu <= _state_ifu_T_1;
    end else begin
      state_ifu <= 2'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_PC = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  state_ifu = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_Cache(
  input         clock,
  input         reset,
  output        from_IFU_ready,
  input         from_IFU_valid,
  input  [31:0] from_IFU_bits_addr,
  output        to_IFU_valid,
  output [31:0] to_IFU_bits_data,
  input         to_sram_ar_ready,
  output        to_sram_ar_valid,
  output [31:0] to_sram_ar_bits_addr,
  output [7:0]  to_sram_ar_bits_len,
  output        to_sram_r_ready,
  input         to_sram_r_valid,
  input  [31:0] to_sram_r_bits_data,
  input         to_sram_r_bits_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2862;
  reg [31:0] _RAND_2865;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2889;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2895;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2943;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2958;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2967;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2973;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3003;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3021;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3045;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3051;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3069;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2905;
  reg [31:0] _RAND_2906;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3055;
  reg [31:0] _RAND_3056;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [31:0] _RAND_3099;
  reg [31:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [31:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [31:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
  reg [31:0] _RAND_3140;
  reg [31:0] _RAND_3141;
  reg [31:0] _RAND_3142;
  reg [31:0] _RAND_3143;
  reg [31:0] _RAND_3144;
  reg [31:0] _RAND_3145;
  reg [31:0] _RAND_3146;
  reg [31:0] _RAND_3147;
  reg [31:0] _RAND_3148;
  reg [31:0] _RAND_3149;
  reg [31:0] _RAND_3150;
  reg [31:0] _RAND_3151;
  reg [31:0] _RAND_3152;
  reg [31:0] _RAND_3153;
  reg [31:0] _RAND_3154;
  reg [31:0] _RAND_3155;
  reg [31:0] _RAND_3156;
  reg [31:0] _RAND_3157;
  reg [31:0] _RAND_3158;
  reg [31:0] _RAND_3159;
  reg [31:0] _RAND_3160;
  reg [31:0] _RAND_3161;
  reg [31:0] _RAND_3162;
  reg [31:0] _RAND_3163;
  reg [31:0] _RAND_3164;
  reg [31:0] _RAND_3165;
  reg [31:0] _RAND_3166;
  reg [31:0] _RAND_3167;
  reg [31:0] _RAND_3168;
  reg [31:0] _RAND_3169;
  reg [31:0] _RAND_3170;
  reg [31:0] _RAND_3171;
  reg [31:0] _RAND_3172;
  reg [31:0] _RAND_3173;
  reg [31:0] _RAND_3174;
  reg [31:0] _RAND_3175;
  reg [31:0] _RAND_3176;
  reg [31:0] _RAND_3177;
  reg [31:0] _RAND_3178;
  reg [31:0] _RAND_3179;
  reg [31:0] _RAND_3180;
  reg [31:0] _RAND_3181;
  reg [31:0] _RAND_3182;
  reg [31:0] _RAND_3183;
  reg [31:0] _RAND_3184;
  reg [31:0] _RAND_3185;
  reg [31:0] _RAND_3186;
  reg [31:0] _RAND_3187;
  reg [31:0] _RAND_3188;
  reg [31:0] _RAND_3189;
  reg [31:0] _RAND_3190;
  reg [31:0] _RAND_3191;
  reg [31:0] _RAND_3192;
  reg [31:0] _RAND_3193;
  reg [31:0] _RAND_3194;
  reg [31:0] _RAND_3195;
  reg [31:0] _RAND_3196;
  reg [31:0] _RAND_3197;
  reg [31:0] _RAND_3198;
  reg [31:0] _RAND_3199;
  reg [31:0] _RAND_3200;
  reg [31:0] _RAND_3201;
  reg [31:0] _RAND_3202;
  reg [31:0] _RAND_3203;
  reg [31:0] _RAND_3204;
  reg [31:0] _RAND_3205;
  reg [31:0] _RAND_3206;
  reg [31:0] _RAND_3207;
  reg [31:0] _RAND_3208;
  reg [31:0] _RAND_3209;
  reg [31:0] _RAND_3210;
  reg [31:0] _RAND_3211;
  reg [31:0] _RAND_3212;
  reg [31:0] _RAND_3213;
  reg [31:0] _RAND_3214;
  reg [31:0] _RAND_3215;
  reg [31:0] _RAND_3216;
  reg [31:0] _RAND_3217;
  reg [31:0] _RAND_3218;
  reg [31:0] _RAND_3219;
  reg [31:0] _RAND_3220;
  reg [31:0] _RAND_3221;
  reg [31:0] _RAND_3222;
  reg [31:0] _RAND_3223;
  reg [31:0] _RAND_3224;
  reg [31:0] _RAND_3225;
  reg [31:0] _RAND_3226;
  reg [31:0] _RAND_3227;
  reg [31:0] _RAND_3228;
  reg [31:0] _RAND_3229;
  reg [31:0] _RAND_3230;
  reg [31:0] _RAND_3231;
  reg [31:0] _RAND_3232;
  reg [31:0] _RAND_3233;
  reg [31:0] _RAND_3234;
  reg [31:0] _RAND_3235;
  reg [31:0] _RAND_3236;
  reg [31:0] _RAND_3237;
  reg [31:0] _RAND_3238;
  reg [31:0] _RAND_3239;
  reg [31:0] _RAND_3240;
  reg [31:0] _RAND_3241;
  reg [31:0] _RAND_3242;
  reg [31:0] _RAND_3243;
  reg [31:0] _RAND_3244;
  reg [31:0] _RAND_3245;
  reg [31:0] _RAND_3246;
  reg [31:0] _RAND_3247;
  reg [31:0] _RAND_3248;
  reg [31:0] _RAND_3249;
  reg [31:0] _RAND_3250;
  reg [31:0] _RAND_3251;
  reg [31:0] _RAND_3252;
  reg [31:0] _RAND_3253;
  reg [31:0] _RAND_3254;
  reg [31:0] _RAND_3255;
  reg [31:0] _RAND_3256;
  reg [31:0] _RAND_3257;
  reg [31:0] _RAND_3258;
  reg [31:0] _RAND_3259;
  reg [31:0] _RAND_3260;
  reg [31:0] _RAND_3261;
  reg [31:0] _RAND_3262;
  reg [31:0] _RAND_3263;
  reg [31:0] _RAND_3264;
  reg [31:0] _RAND_3265;
  reg [31:0] _RAND_3266;
  reg [31:0] _RAND_3267;
  reg [31:0] _RAND_3268;
  reg [31:0] _RAND_3269;
  reg [31:0] _RAND_3270;
  reg [31:0] _RAND_3271;
  reg [31:0] _RAND_3272;
  reg [31:0] _RAND_3273;
  reg [31:0] _RAND_3274;
  reg [31:0] _RAND_3275;
  reg [31:0] _RAND_3276;
  reg [31:0] _RAND_3277;
  reg [31:0] _RAND_3278;
  reg [31:0] _RAND_3279;
  reg [31:0] _RAND_3280;
  reg [31:0] _RAND_3281;
  reg [31:0] _RAND_3282;
  reg [31:0] _RAND_3283;
  reg [31:0] _RAND_3284;
  reg [31:0] _RAND_3285;
  reg [31:0] _RAND_3286;
  reg [31:0] _RAND_3287;
  reg [31:0] _RAND_3288;
  reg [31:0] _RAND_3289;
  reg [31:0] _RAND_3290;
  reg [31:0] _RAND_3291;
  reg [31:0] _RAND_3292;
  reg [31:0] _RAND_3293;
  reg [31:0] _RAND_3294;
  reg [31:0] _RAND_3295;
  reg [31:0] _RAND_3296;
  reg [31:0] _RAND_3297;
  reg [31:0] _RAND_3298;
  reg [31:0] _RAND_3299;
  reg [31:0] _RAND_3300;
  reg [31:0] _RAND_3301;
  reg [31:0] _RAND_3302;
  reg [31:0] _RAND_3303;
  reg [31:0] _RAND_3304;
  reg [31:0] _RAND_3305;
  reg [31:0] _RAND_3306;
  reg [31:0] _RAND_3307;
  reg [31:0] _RAND_3308;
  reg [31:0] _RAND_3309;
  reg [31:0] _RAND_3310;
  reg [31:0] _RAND_3311;
  reg [31:0] _RAND_3312;
  reg [31:0] _RAND_3313;
  reg [31:0] _RAND_3314;
  reg [31:0] _RAND_3315;
  reg [31:0] _RAND_3316;
  reg [31:0] _RAND_3317;
  reg [31:0] _RAND_3318;
  reg [31:0] _RAND_3319;
  reg [31:0] _RAND_3320;
  reg [31:0] _RAND_3321;
  reg [31:0] _RAND_3322;
  reg [31:0] _RAND_3323;
  reg [31:0] _RAND_3324;
  reg [31:0] _RAND_3325;
  reg [31:0] _RAND_3326;
  reg [31:0] _RAND_3327;
  reg [31:0] _RAND_3328;
  reg [31:0] _RAND_3329;
  reg [31:0] _RAND_3330;
  reg [31:0] _RAND_3331;
  reg [31:0] _RAND_3332;
  reg [31:0] _RAND_3333;
  reg [31:0] _RAND_3334;
  reg [31:0] _RAND_3335;
  reg [31:0] _RAND_3336;
  reg [31:0] _RAND_3337;
  reg [31:0] _RAND_3338;
  reg [31:0] _RAND_3339;
  reg [31:0] _RAND_3340;
  reg [31:0] _RAND_3341;
  reg [31:0] _RAND_3342;
  reg [31:0] _RAND_3343;
  reg [31:0] _RAND_3344;
  reg [31:0] _RAND_3345;
  reg [31:0] _RAND_3346;
  reg [31:0] _RAND_3347;
  reg [31:0] _RAND_3348;
  reg [31:0] _RAND_3349;
  reg [31:0] _RAND_3350;
  reg [31:0] _RAND_3351;
  reg [31:0] _RAND_3352;
  reg [31:0] _RAND_3353;
  reg [31:0] _RAND_3354;
  reg [31:0] _RAND_3355;
  reg [31:0] _RAND_3356;
  reg [31:0] _RAND_3357;
  reg [31:0] _RAND_3358;
  reg [31:0] _RAND_3359;
  reg [31:0] _RAND_3360;
  reg [31:0] _RAND_3361;
  reg [31:0] _RAND_3362;
  reg [31:0] _RAND_3363;
  reg [31:0] _RAND_3364;
  reg [31:0] _RAND_3365;
  reg [31:0] _RAND_3366;
  reg [31:0] _RAND_3367;
  reg [31:0] _RAND_3368;
  reg [31:0] _RAND_3369;
  reg [31:0] _RAND_3370;
  reg [31:0] _RAND_3371;
  reg [31:0] _RAND_3372;
  reg [31:0] _RAND_3373;
  reg [31:0] _RAND_3374;
  reg [31:0] _RAND_3375;
  reg [31:0] _RAND_3376;
  reg [31:0] _RAND_3377;
  reg [31:0] _RAND_3378;
  reg [31:0] _RAND_3379;
  reg [31:0] _RAND_3380;
  reg [31:0] _RAND_3381;
  reg [31:0] _RAND_3382;
  reg [31:0] _RAND_3383;
  reg [31:0] _RAND_3384;
  reg [31:0] _RAND_3385;
  reg [31:0] _RAND_3386;
  reg [31:0] _RAND_3387;
  reg [31:0] _RAND_3388;
  reg [31:0] _RAND_3389;
  reg [31:0] _RAND_3390;
  reg [31:0] _RAND_3391;
  reg [31:0] _RAND_3392;
  reg [31:0] _RAND_3393;
  reg [31:0] _RAND_3394;
  reg [31:0] _RAND_3395;
  reg [31:0] _RAND_3396;
  reg [31:0] _RAND_3397;
  reg [31:0] _RAND_3398;
  reg [31:0] _RAND_3399;
  reg [31:0] _RAND_3400;
  reg [31:0] _RAND_3401;
  reg [31:0] _RAND_3402;
  reg [31:0] _RAND_3403;
  reg [31:0] _RAND_3404;
  reg [31:0] _RAND_3405;
  reg [31:0] _RAND_3406;
  reg [31:0] _RAND_3407;
  reg [31:0] _RAND_3408;
  reg [31:0] _RAND_3409;
  reg [31:0] _RAND_3410;
  reg [31:0] _RAND_3411;
  reg [31:0] _RAND_3412;
  reg [31:0] _RAND_3413;
  reg [31:0] _RAND_3414;
  reg [31:0] _RAND_3415;
  reg [31:0] _RAND_3416;
  reg [31:0] _RAND_3417;
  reg [31:0] _RAND_3418;
  reg [31:0] _RAND_3419;
  reg [31:0] _RAND_3420;
  reg [31:0] _RAND_3421;
  reg [31:0] _RAND_3422;
  reg [31:0] _RAND_3423;
  reg [31:0] _RAND_3424;
  reg [31:0] _RAND_3425;
  reg [31:0] _RAND_3426;
  reg [31:0] _RAND_3427;
  reg [31:0] _RAND_3428;
  reg [31:0] _RAND_3429;
  reg [31:0] _RAND_3430;
  reg [31:0] _RAND_3431;
  reg [31:0] _RAND_3432;
  reg [31:0] _RAND_3433;
  reg [31:0] _RAND_3434;
  reg [31:0] _RAND_3435;
  reg [31:0] _RAND_3436;
  reg [31:0] _RAND_3437;
  reg [31:0] _RAND_3438;
  reg [31:0] _RAND_3439;
  reg [31:0] _RAND_3440;
  reg [31:0] _RAND_3441;
  reg [31:0] _RAND_3442;
  reg [31:0] _RAND_3443;
  reg [31:0] _RAND_3444;
  reg [31:0] _RAND_3445;
  reg [31:0] _RAND_3446;
  reg [31:0] _RAND_3447;
  reg [31:0] _RAND_3448;
  reg [31:0] _RAND_3449;
  reg [31:0] _RAND_3450;
  reg [31:0] _RAND_3451;
  reg [31:0] _RAND_3452;
  reg [31:0] _RAND_3453;
  reg [31:0] _RAND_3454;
  reg [31:0] _RAND_3455;
  reg [31:0] _RAND_3456;
  reg [31:0] _RAND_3457;
  reg [31:0] _RAND_3458;
  reg [31:0] _RAND_3459;
  reg [31:0] _RAND_3460;
  reg [31:0] _RAND_3461;
  reg [31:0] _RAND_3462;
  reg [31:0] _RAND_3463;
  reg [31:0] _RAND_3464;
  reg [31:0] _RAND_3465;
  reg [31:0] _RAND_3466;
  reg [31:0] _RAND_3467;
  reg [31:0] _RAND_3468;
  reg [31:0] _RAND_3469;
  reg [31:0] _RAND_3470;
  reg [31:0] _RAND_3471;
  reg [31:0] _RAND_3472;
  reg [31:0] _RAND_3473;
  reg [31:0] _RAND_3474;
  reg [31:0] _RAND_3475;
  reg [31:0] _RAND_3476;
  reg [31:0] _RAND_3477;
  reg [31:0] _RAND_3478;
  reg [31:0] _RAND_3479;
  reg [31:0] _RAND_3480;
  reg [31:0] _RAND_3481;
  reg [31:0] _RAND_3482;
  reg [31:0] _RAND_3483;
  reg [31:0] _RAND_3484;
  reg [31:0] _RAND_3485;
  reg [31:0] _RAND_3486;
  reg [31:0] _RAND_3487;
  reg [31:0] _RAND_3488;
  reg [31:0] _RAND_3489;
  reg [31:0] _RAND_3490;
  reg [31:0] _RAND_3491;
  reg [31:0] _RAND_3492;
  reg [31:0] _RAND_3493;
  reg [31:0] _RAND_3494;
  reg [31:0] _RAND_3495;
  reg [31:0] _RAND_3496;
  reg [31:0] _RAND_3497;
  reg [31:0] _RAND_3498;
  reg [31:0] _RAND_3499;
  reg [31:0] _RAND_3500;
  reg [31:0] _RAND_3501;
  reg [31:0] _RAND_3502;
  reg [31:0] _RAND_3503;
  reg [31:0] _RAND_3504;
  reg [31:0] _RAND_3505;
  reg [31:0] _RAND_3506;
  reg [31:0] _RAND_3507;
  reg [31:0] _RAND_3508;
  reg [31:0] _RAND_3509;
  reg [31:0] _RAND_3510;
  reg [31:0] _RAND_3511;
  reg [31:0] _RAND_3512;
  reg [31:0] _RAND_3513;
  reg [31:0] _RAND_3514;
  reg [31:0] _RAND_3515;
  reg [31:0] _RAND_3516;
  reg [31:0] _RAND_3517;
  reg [31:0] _RAND_3518;
  reg [31:0] _RAND_3519;
  reg [31:0] _RAND_3520;
  reg [31:0] _RAND_3521;
  reg [31:0] _RAND_3522;
  reg [31:0] _RAND_3523;
  reg [31:0] _RAND_3524;
  reg [31:0] _RAND_3525;
  reg [31:0] _RAND_3526;
  reg [31:0] _RAND_3527;
  reg [31:0] _RAND_3528;
  reg [31:0] _RAND_3529;
  reg [31:0] _RAND_3530;
  reg [31:0] _RAND_3531;
  reg [31:0] _RAND_3532;
  reg [31:0] _RAND_3533;
  reg [31:0] _RAND_3534;
  reg [31:0] _RAND_3535;
  reg [31:0] _RAND_3536;
  reg [31:0] _RAND_3537;
  reg [31:0] _RAND_3538;
  reg [31:0] _RAND_3539;
  reg [31:0] _RAND_3540;
  reg [31:0] _RAND_3541;
  reg [31:0] _RAND_3542;
  reg [31:0] _RAND_3543;
  reg [31:0] _RAND_3544;
  reg [31:0] _RAND_3545;
  reg [31:0] _RAND_3546;
  reg [31:0] _RAND_3547;
  reg [31:0] _RAND_3548;
  reg [31:0] _RAND_3549;
  reg [31:0] _RAND_3550;
  reg [31:0] _RAND_3551;
  reg [31:0] _RAND_3552;
  reg [31:0] _RAND_3553;
  reg [31:0] _RAND_3554;
  reg [31:0] _RAND_3555;
  reg [31:0] _RAND_3556;
  reg [31:0] _RAND_3557;
  reg [31:0] _RAND_3558;
  reg [31:0] _RAND_3559;
  reg [31:0] _RAND_3560;
  reg [31:0] _RAND_3561;
  reg [31:0] _RAND_3562;
  reg [31:0] _RAND_3563;
  reg [31:0] _RAND_3564;
  reg [31:0] _RAND_3565;
  reg [31:0] _RAND_3566;
  reg [31:0] _RAND_3567;
  reg [31:0] _RAND_3568;
  reg [31:0] _RAND_3569;
  reg [31:0] _RAND_3570;
  reg [31:0] _RAND_3571;
  reg [31:0] _RAND_3572;
  reg [31:0] _RAND_3573;
  reg [31:0] _RAND_3574;
  reg [31:0] _RAND_3575;
  reg [31:0] _RAND_3576;
  reg [31:0] _RAND_3577;
  reg [31:0] _RAND_3578;
  reg [31:0] _RAND_3579;
  reg [31:0] _RAND_3580;
  reg [31:0] _RAND_3581;
  reg [31:0] _RAND_3582;
  reg [31:0] _RAND_3583;
  reg [31:0] _RAND_3584;
  reg [31:0] _RAND_3585;
  reg [31:0] _RAND_3586;
  reg [31:0] _RAND_3587;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] dataArray_0_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_0_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_0_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_0_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_1_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_1_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_1_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_2_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_2_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_2_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_3_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_3_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_3_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_4_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_4_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_4_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_5_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_5_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_5_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_6_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_6_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_6_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_7_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_7_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_7_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_8_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_8_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_8_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_9_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_9_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_9_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_10_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_10_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_10_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_11_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_11_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_11_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_12_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_12_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_12_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_13_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_13_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_13_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_14_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_14_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_14_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_15_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_15_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_15_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_16_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_16_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_16_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_16_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_16_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_16_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_16_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_16_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_17_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_17_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_17_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_17_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_17_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_17_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_17_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_17_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_18_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_18_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_18_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_18_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_18_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_18_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_18_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_18_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_19_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_19_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_19_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_19_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_19_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_19_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_19_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_19_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_20_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_20_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_20_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_20_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_20_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_20_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_20_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_20_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_21_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_21_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_21_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_21_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_21_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_21_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_21_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_21_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_22_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_22_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_22_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_22_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_22_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_22_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_22_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_22_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_23_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_23_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_23_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_23_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_23_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_23_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_23_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_23_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_24_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_24_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_24_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_24_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_24_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_24_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_24_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_24_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_25_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_25_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_25_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_25_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_25_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_25_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_25_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_25_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_26_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_26_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_26_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_26_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_26_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_26_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_26_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_26_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_27_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_27_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_27_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_27_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_27_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_27_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_27_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_27_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_28_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_28_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_28_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_28_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_28_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_28_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_28_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_28_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_29_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_29_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_29_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_29_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_29_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_29_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_29_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_29_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_30_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_30_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_30_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_30_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_30_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_30_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_30_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_30_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_31_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_31_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_31_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_31_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_31_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_31_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_31_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_31_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_32_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_32_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_32_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_32_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_32_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_32_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_32_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_32_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_33_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_33_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_33_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_33_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_33_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_33_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_33_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_33_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_34_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_34_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_34_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_34_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_34_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_34_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_34_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_34_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_35_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_35_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_35_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_35_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_35_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_35_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_35_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_35_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_36_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_36_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_36_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_36_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_36_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_36_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_36_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_36_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_37_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_37_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_37_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_37_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_37_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_37_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_37_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_37_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_38_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_38_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_38_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_38_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_38_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_38_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_38_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_38_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_39_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_39_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_39_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_39_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_39_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_39_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_39_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_39_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_40_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_40_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_40_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_40_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_40_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_40_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_40_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_40_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_41_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_41_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_41_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_41_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_41_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_41_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_41_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_41_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_42_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_42_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_42_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_42_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_42_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_42_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_42_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_42_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_43_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_43_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_43_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_43_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_43_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_43_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_43_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_43_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_44_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_44_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_44_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_44_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_44_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_44_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_44_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_44_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_45_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_45_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_45_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_45_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_45_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_45_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_45_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_45_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_46_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_46_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_46_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_46_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_46_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_46_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_46_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_46_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_47_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_47_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_47_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_47_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_47_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_47_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_47_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_47_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_48_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_48_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_48_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_48_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_48_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_48_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_48_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_48_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_49_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_49_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_49_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_49_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_49_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_49_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_49_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_49_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_50_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_50_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_50_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_50_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_50_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_50_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_50_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_50_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_51_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_51_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_51_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_51_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_51_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_51_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_51_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_51_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_52_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_52_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_52_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_52_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_52_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_52_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_52_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_52_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_53_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_53_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_53_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_53_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_53_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_53_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_53_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_53_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_54_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_54_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_54_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_54_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_54_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_54_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_54_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_54_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_55_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_55_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_55_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_55_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_55_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_55_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_55_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_55_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_56_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_56_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_56_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_56_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_56_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_56_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_56_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_56_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_57_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_57_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_57_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_57_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_57_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_57_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_57_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_57_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_58_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_58_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_58_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_58_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_58_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_58_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_58_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_58_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_59_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_59_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_59_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_59_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_59_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_59_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_59_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_59_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_60_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_60_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_60_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_60_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_60_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_60_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_60_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_60_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_61_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_61_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_61_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_61_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_61_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_61_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_61_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_61_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_62_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_62_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_62_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_62_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_62_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_62_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_62_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_62_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_0 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_0_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_0_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_1 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_1_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_1_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_2 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_2_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_2_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_3 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_3_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_3_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_4 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_4_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_4_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_5 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_5_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_5_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_6 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_6_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_6_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_7 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_7_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_7_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_8 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_8_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_8_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_9 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_9_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_9_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_10 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_10_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_10_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_11 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_11_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_11_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_12 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_12_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_12_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_13 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_13_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_13_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_14 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_14_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_14_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_63_15 [0:3]; // @[cache.scala 30:33]
  wire  dataArray_63_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_63_15_MPORT_data; // @[cache.scala 30:33]
  wire [1:0] dataArray_63_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_63_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_63_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_63_15_cachedata_MPORT_en_pipe_0;
  reg [1:0] dataArray_63_15_cachedata_MPORT_addr_pipe_0;
  reg [1:0] replace_set; // @[cache.scala 21:30]
  wire [5:0] EntId = from_IFU_bits_addr[5:0] / 3'h4; // @[cache.scala 22:59]
  wire [5:0] CacheLineId = from_IFU_bits_addr[11:6]; // @[cache.scala 23:41]
  wire [19:0] tag = from_IFU_bits_addr[31:12]; // @[cache.scala 24:39]
  reg [1:0] random_num; // @[cache.scala 27:29]
  wire [1:0] _random_num_T_1 = random_num + 2'h1; // @[cache.scala 28:29]
  reg [19:0] tagArray_0_0; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_1; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_2; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_3; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_4; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_5; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_6; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_7; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_8; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_9; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_10; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_11; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_12; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_13; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_14; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_15; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_16; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_17; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_18; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_19; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_20; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_21; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_22; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_23; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_24; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_25; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_26; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_27; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_28; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_29; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_30; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_31; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_32; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_33; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_34; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_35; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_36; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_37; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_38; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_39; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_40; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_41; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_42; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_43; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_44; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_45; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_46; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_47; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_48; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_49; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_50; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_51; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_52; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_53; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_54; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_55; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_56; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_57; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_58; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_59; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_60; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_61; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_62; // @[cache.scala 31:29]
  reg [19:0] tagArray_0_63; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_0; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_1; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_2; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_3; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_4; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_5; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_6; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_7; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_8; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_9; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_10; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_11; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_12; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_13; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_14; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_15; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_16; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_17; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_18; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_19; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_20; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_21; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_22; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_23; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_24; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_25; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_26; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_27; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_28; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_29; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_30; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_31; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_32; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_33; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_34; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_35; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_36; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_37; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_38; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_39; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_40; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_41; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_42; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_43; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_44; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_45; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_46; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_47; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_48; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_49; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_50; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_51; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_52; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_53; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_54; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_55; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_56; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_57; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_58; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_59; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_60; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_61; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_62; // @[cache.scala 31:29]
  reg [19:0] tagArray_1_63; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_0; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_1; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_2; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_3; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_4; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_5; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_6; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_7; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_8; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_9; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_10; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_11; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_12; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_13; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_14; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_15; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_16; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_17; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_18; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_19; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_20; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_21; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_22; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_23; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_24; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_25; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_26; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_27; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_28; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_29; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_30; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_31; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_32; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_33; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_34; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_35; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_36; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_37; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_38; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_39; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_40; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_41; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_42; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_43; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_44; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_45; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_46; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_47; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_48; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_49; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_50; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_51; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_52; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_53; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_54; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_55; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_56; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_57; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_58; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_59; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_60; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_61; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_62; // @[cache.scala 31:29]
  reg [19:0] tagArray_2_63; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_0; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_1; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_2; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_3; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_4; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_5; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_6; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_7; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_8; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_9; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_10; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_11; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_12; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_13; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_14; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_15; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_16; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_17; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_18; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_19; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_20; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_21; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_22; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_23; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_24; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_25; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_26; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_27; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_28; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_29; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_30; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_31; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_32; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_33; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_34; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_35; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_36; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_37; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_38; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_39; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_40; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_41; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_42; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_43; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_44; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_45; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_46; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_47; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_48; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_49; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_50; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_51; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_52; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_53; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_54; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_55; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_56; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_57; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_58; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_59; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_60; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_61; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_62; // @[cache.scala 31:29]
  reg [19:0] tagArray_3_63; // @[cache.scala 31:29]
  reg  validArray_0_0; // @[cache.scala 32:29]
  reg  validArray_0_1; // @[cache.scala 32:29]
  reg  validArray_0_2; // @[cache.scala 32:29]
  reg  validArray_0_3; // @[cache.scala 32:29]
  reg  validArray_0_4; // @[cache.scala 32:29]
  reg  validArray_0_5; // @[cache.scala 32:29]
  reg  validArray_0_6; // @[cache.scala 32:29]
  reg  validArray_0_7; // @[cache.scala 32:29]
  reg  validArray_0_8; // @[cache.scala 32:29]
  reg  validArray_0_9; // @[cache.scala 32:29]
  reg  validArray_0_10; // @[cache.scala 32:29]
  reg  validArray_0_11; // @[cache.scala 32:29]
  reg  validArray_0_12; // @[cache.scala 32:29]
  reg  validArray_0_13; // @[cache.scala 32:29]
  reg  validArray_0_14; // @[cache.scala 32:29]
  reg  validArray_0_15; // @[cache.scala 32:29]
  reg  validArray_0_16; // @[cache.scala 32:29]
  reg  validArray_0_17; // @[cache.scala 32:29]
  reg  validArray_0_18; // @[cache.scala 32:29]
  reg  validArray_0_19; // @[cache.scala 32:29]
  reg  validArray_0_20; // @[cache.scala 32:29]
  reg  validArray_0_21; // @[cache.scala 32:29]
  reg  validArray_0_22; // @[cache.scala 32:29]
  reg  validArray_0_23; // @[cache.scala 32:29]
  reg  validArray_0_24; // @[cache.scala 32:29]
  reg  validArray_0_25; // @[cache.scala 32:29]
  reg  validArray_0_26; // @[cache.scala 32:29]
  reg  validArray_0_27; // @[cache.scala 32:29]
  reg  validArray_0_28; // @[cache.scala 32:29]
  reg  validArray_0_29; // @[cache.scala 32:29]
  reg  validArray_0_30; // @[cache.scala 32:29]
  reg  validArray_0_31; // @[cache.scala 32:29]
  reg  validArray_0_32; // @[cache.scala 32:29]
  reg  validArray_0_33; // @[cache.scala 32:29]
  reg  validArray_0_34; // @[cache.scala 32:29]
  reg  validArray_0_35; // @[cache.scala 32:29]
  reg  validArray_0_36; // @[cache.scala 32:29]
  reg  validArray_0_37; // @[cache.scala 32:29]
  reg  validArray_0_38; // @[cache.scala 32:29]
  reg  validArray_0_39; // @[cache.scala 32:29]
  reg  validArray_0_40; // @[cache.scala 32:29]
  reg  validArray_0_41; // @[cache.scala 32:29]
  reg  validArray_0_42; // @[cache.scala 32:29]
  reg  validArray_0_43; // @[cache.scala 32:29]
  reg  validArray_0_44; // @[cache.scala 32:29]
  reg  validArray_0_45; // @[cache.scala 32:29]
  reg  validArray_0_46; // @[cache.scala 32:29]
  reg  validArray_0_47; // @[cache.scala 32:29]
  reg  validArray_0_48; // @[cache.scala 32:29]
  reg  validArray_0_49; // @[cache.scala 32:29]
  reg  validArray_0_50; // @[cache.scala 32:29]
  reg  validArray_0_51; // @[cache.scala 32:29]
  reg  validArray_0_52; // @[cache.scala 32:29]
  reg  validArray_0_53; // @[cache.scala 32:29]
  reg  validArray_0_54; // @[cache.scala 32:29]
  reg  validArray_0_55; // @[cache.scala 32:29]
  reg  validArray_0_56; // @[cache.scala 32:29]
  reg  validArray_0_57; // @[cache.scala 32:29]
  reg  validArray_0_58; // @[cache.scala 32:29]
  reg  validArray_0_59; // @[cache.scala 32:29]
  reg  validArray_0_60; // @[cache.scala 32:29]
  reg  validArray_0_61; // @[cache.scala 32:29]
  reg  validArray_0_62; // @[cache.scala 32:29]
  reg  validArray_0_63; // @[cache.scala 32:29]
  reg  validArray_1_0; // @[cache.scala 32:29]
  reg  validArray_1_1; // @[cache.scala 32:29]
  reg  validArray_1_2; // @[cache.scala 32:29]
  reg  validArray_1_3; // @[cache.scala 32:29]
  reg  validArray_1_4; // @[cache.scala 32:29]
  reg  validArray_1_5; // @[cache.scala 32:29]
  reg  validArray_1_6; // @[cache.scala 32:29]
  reg  validArray_1_7; // @[cache.scala 32:29]
  reg  validArray_1_8; // @[cache.scala 32:29]
  reg  validArray_1_9; // @[cache.scala 32:29]
  reg  validArray_1_10; // @[cache.scala 32:29]
  reg  validArray_1_11; // @[cache.scala 32:29]
  reg  validArray_1_12; // @[cache.scala 32:29]
  reg  validArray_1_13; // @[cache.scala 32:29]
  reg  validArray_1_14; // @[cache.scala 32:29]
  reg  validArray_1_15; // @[cache.scala 32:29]
  reg  validArray_1_16; // @[cache.scala 32:29]
  reg  validArray_1_17; // @[cache.scala 32:29]
  reg  validArray_1_18; // @[cache.scala 32:29]
  reg  validArray_1_19; // @[cache.scala 32:29]
  reg  validArray_1_20; // @[cache.scala 32:29]
  reg  validArray_1_21; // @[cache.scala 32:29]
  reg  validArray_1_22; // @[cache.scala 32:29]
  reg  validArray_1_23; // @[cache.scala 32:29]
  reg  validArray_1_24; // @[cache.scala 32:29]
  reg  validArray_1_25; // @[cache.scala 32:29]
  reg  validArray_1_26; // @[cache.scala 32:29]
  reg  validArray_1_27; // @[cache.scala 32:29]
  reg  validArray_1_28; // @[cache.scala 32:29]
  reg  validArray_1_29; // @[cache.scala 32:29]
  reg  validArray_1_30; // @[cache.scala 32:29]
  reg  validArray_1_31; // @[cache.scala 32:29]
  reg  validArray_1_32; // @[cache.scala 32:29]
  reg  validArray_1_33; // @[cache.scala 32:29]
  reg  validArray_1_34; // @[cache.scala 32:29]
  reg  validArray_1_35; // @[cache.scala 32:29]
  reg  validArray_1_36; // @[cache.scala 32:29]
  reg  validArray_1_37; // @[cache.scala 32:29]
  reg  validArray_1_38; // @[cache.scala 32:29]
  reg  validArray_1_39; // @[cache.scala 32:29]
  reg  validArray_1_40; // @[cache.scala 32:29]
  reg  validArray_1_41; // @[cache.scala 32:29]
  reg  validArray_1_42; // @[cache.scala 32:29]
  reg  validArray_1_43; // @[cache.scala 32:29]
  reg  validArray_1_44; // @[cache.scala 32:29]
  reg  validArray_1_45; // @[cache.scala 32:29]
  reg  validArray_1_46; // @[cache.scala 32:29]
  reg  validArray_1_47; // @[cache.scala 32:29]
  reg  validArray_1_48; // @[cache.scala 32:29]
  reg  validArray_1_49; // @[cache.scala 32:29]
  reg  validArray_1_50; // @[cache.scala 32:29]
  reg  validArray_1_51; // @[cache.scala 32:29]
  reg  validArray_1_52; // @[cache.scala 32:29]
  reg  validArray_1_53; // @[cache.scala 32:29]
  reg  validArray_1_54; // @[cache.scala 32:29]
  reg  validArray_1_55; // @[cache.scala 32:29]
  reg  validArray_1_56; // @[cache.scala 32:29]
  reg  validArray_1_57; // @[cache.scala 32:29]
  reg  validArray_1_58; // @[cache.scala 32:29]
  reg  validArray_1_59; // @[cache.scala 32:29]
  reg  validArray_1_60; // @[cache.scala 32:29]
  reg  validArray_1_61; // @[cache.scala 32:29]
  reg  validArray_1_62; // @[cache.scala 32:29]
  reg  validArray_1_63; // @[cache.scala 32:29]
  reg  validArray_2_0; // @[cache.scala 32:29]
  reg  validArray_2_1; // @[cache.scala 32:29]
  reg  validArray_2_2; // @[cache.scala 32:29]
  reg  validArray_2_3; // @[cache.scala 32:29]
  reg  validArray_2_4; // @[cache.scala 32:29]
  reg  validArray_2_5; // @[cache.scala 32:29]
  reg  validArray_2_6; // @[cache.scala 32:29]
  reg  validArray_2_7; // @[cache.scala 32:29]
  reg  validArray_2_8; // @[cache.scala 32:29]
  reg  validArray_2_9; // @[cache.scala 32:29]
  reg  validArray_2_10; // @[cache.scala 32:29]
  reg  validArray_2_11; // @[cache.scala 32:29]
  reg  validArray_2_12; // @[cache.scala 32:29]
  reg  validArray_2_13; // @[cache.scala 32:29]
  reg  validArray_2_14; // @[cache.scala 32:29]
  reg  validArray_2_15; // @[cache.scala 32:29]
  reg  validArray_2_16; // @[cache.scala 32:29]
  reg  validArray_2_17; // @[cache.scala 32:29]
  reg  validArray_2_18; // @[cache.scala 32:29]
  reg  validArray_2_19; // @[cache.scala 32:29]
  reg  validArray_2_20; // @[cache.scala 32:29]
  reg  validArray_2_21; // @[cache.scala 32:29]
  reg  validArray_2_22; // @[cache.scala 32:29]
  reg  validArray_2_23; // @[cache.scala 32:29]
  reg  validArray_2_24; // @[cache.scala 32:29]
  reg  validArray_2_25; // @[cache.scala 32:29]
  reg  validArray_2_26; // @[cache.scala 32:29]
  reg  validArray_2_27; // @[cache.scala 32:29]
  reg  validArray_2_28; // @[cache.scala 32:29]
  reg  validArray_2_29; // @[cache.scala 32:29]
  reg  validArray_2_30; // @[cache.scala 32:29]
  reg  validArray_2_31; // @[cache.scala 32:29]
  reg  validArray_2_32; // @[cache.scala 32:29]
  reg  validArray_2_33; // @[cache.scala 32:29]
  reg  validArray_2_34; // @[cache.scala 32:29]
  reg  validArray_2_35; // @[cache.scala 32:29]
  reg  validArray_2_36; // @[cache.scala 32:29]
  reg  validArray_2_37; // @[cache.scala 32:29]
  reg  validArray_2_38; // @[cache.scala 32:29]
  reg  validArray_2_39; // @[cache.scala 32:29]
  reg  validArray_2_40; // @[cache.scala 32:29]
  reg  validArray_2_41; // @[cache.scala 32:29]
  reg  validArray_2_42; // @[cache.scala 32:29]
  reg  validArray_2_43; // @[cache.scala 32:29]
  reg  validArray_2_44; // @[cache.scala 32:29]
  reg  validArray_2_45; // @[cache.scala 32:29]
  reg  validArray_2_46; // @[cache.scala 32:29]
  reg  validArray_2_47; // @[cache.scala 32:29]
  reg  validArray_2_48; // @[cache.scala 32:29]
  reg  validArray_2_49; // @[cache.scala 32:29]
  reg  validArray_2_50; // @[cache.scala 32:29]
  reg  validArray_2_51; // @[cache.scala 32:29]
  reg  validArray_2_52; // @[cache.scala 32:29]
  reg  validArray_2_53; // @[cache.scala 32:29]
  reg  validArray_2_54; // @[cache.scala 32:29]
  reg  validArray_2_55; // @[cache.scala 32:29]
  reg  validArray_2_56; // @[cache.scala 32:29]
  reg  validArray_2_57; // @[cache.scala 32:29]
  reg  validArray_2_58; // @[cache.scala 32:29]
  reg  validArray_2_59; // @[cache.scala 32:29]
  reg  validArray_2_60; // @[cache.scala 32:29]
  reg  validArray_2_61; // @[cache.scala 32:29]
  reg  validArray_2_62; // @[cache.scala 32:29]
  reg  validArray_2_63; // @[cache.scala 32:29]
  reg  validArray_3_0; // @[cache.scala 32:29]
  reg  validArray_3_1; // @[cache.scala 32:29]
  reg  validArray_3_2; // @[cache.scala 32:29]
  reg  validArray_3_3; // @[cache.scala 32:29]
  reg  validArray_3_4; // @[cache.scala 32:29]
  reg  validArray_3_5; // @[cache.scala 32:29]
  reg  validArray_3_6; // @[cache.scala 32:29]
  reg  validArray_3_7; // @[cache.scala 32:29]
  reg  validArray_3_8; // @[cache.scala 32:29]
  reg  validArray_3_9; // @[cache.scala 32:29]
  reg  validArray_3_10; // @[cache.scala 32:29]
  reg  validArray_3_11; // @[cache.scala 32:29]
  reg  validArray_3_12; // @[cache.scala 32:29]
  reg  validArray_3_13; // @[cache.scala 32:29]
  reg  validArray_3_14; // @[cache.scala 32:29]
  reg  validArray_3_15; // @[cache.scala 32:29]
  reg  validArray_3_16; // @[cache.scala 32:29]
  reg  validArray_3_17; // @[cache.scala 32:29]
  reg  validArray_3_18; // @[cache.scala 32:29]
  reg  validArray_3_19; // @[cache.scala 32:29]
  reg  validArray_3_20; // @[cache.scala 32:29]
  reg  validArray_3_21; // @[cache.scala 32:29]
  reg  validArray_3_22; // @[cache.scala 32:29]
  reg  validArray_3_23; // @[cache.scala 32:29]
  reg  validArray_3_24; // @[cache.scala 32:29]
  reg  validArray_3_25; // @[cache.scala 32:29]
  reg  validArray_3_26; // @[cache.scala 32:29]
  reg  validArray_3_27; // @[cache.scala 32:29]
  reg  validArray_3_28; // @[cache.scala 32:29]
  reg  validArray_3_29; // @[cache.scala 32:29]
  reg  validArray_3_30; // @[cache.scala 32:29]
  reg  validArray_3_31; // @[cache.scala 32:29]
  reg  validArray_3_32; // @[cache.scala 32:29]
  reg  validArray_3_33; // @[cache.scala 32:29]
  reg  validArray_3_34; // @[cache.scala 32:29]
  reg  validArray_3_35; // @[cache.scala 32:29]
  reg  validArray_3_36; // @[cache.scala 32:29]
  reg  validArray_3_37; // @[cache.scala 32:29]
  reg  validArray_3_38; // @[cache.scala 32:29]
  reg  validArray_3_39; // @[cache.scala 32:29]
  reg  validArray_3_40; // @[cache.scala 32:29]
  reg  validArray_3_41; // @[cache.scala 32:29]
  reg  validArray_3_42; // @[cache.scala 32:29]
  reg  validArray_3_43; // @[cache.scala 32:29]
  reg  validArray_3_44; // @[cache.scala 32:29]
  reg  validArray_3_45; // @[cache.scala 32:29]
  reg  validArray_3_46; // @[cache.scala 32:29]
  reg  validArray_3_47; // @[cache.scala 32:29]
  reg  validArray_3_48; // @[cache.scala 32:29]
  reg  validArray_3_49; // @[cache.scala 32:29]
  reg  validArray_3_50; // @[cache.scala 32:29]
  reg  validArray_3_51; // @[cache.scala 32:29]
  reg  validArray_3_52; // @[cache.scala 32:29]
  reg  validArray_3_53; // @[cache.scala 32:29]
  reg  validArray_3_54; // @[cache.scala 32:29]
  reg  validArray_3_55; // @[cache.scala 32:29]
  reg  validArray_3_56; // @[cache.scala 32:29]
  reg  validArray_3_57; // @[cache.scala 32:29]
  reg  validArray_3_58; // @[cache.scala 32:29]
  reg  validArray_3_59; // @[cache.scala 32:29]
  reg  validArray_3_60; // @[cache.scala 32:29]
  reg  validArray_3_61; // @[cache.scala 32:29]
  reg  validArray_3_62; // @[cache.scala 32:29]
  reg  validArray_3_63; // @[cache.scala 32:29]
  wire [19:0] _GEN_1 = 6'h1 == CacheLineId ? tagArray_0_1 : tagArray_0_0; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_2 = 6'h2 == CacheLineId ? tagArray_0_2 : _GEN_1; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_3 = 6'h3 == CacheLineId ? tagArray_0_3 : _GEN_2; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_4 = 6'h4 == CacheLineId ? tagArray_0_4 : _GEN_3; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_5 = 6'h5 == CacheLineId ? tagArray_0_5 : _GEN_4; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_6 = 6'h6 == CacheLineId ? tagArray_0_6 : _GEN_5; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_7 = 6'h7 == CacheLineId ? tagArray_0_7 : _GEN_6; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_8 = 6'h8 == CacheLineId ? tagArray_0_8 : _GEN_7; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_9 = 6'h9 == CacheLineId ? tagArray_0_9 : _GEN_8; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_10 = 6'ha == CacheLineId ? tagArray_0_10 : _GEN_9; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_11 = 6'hb == CacheLineId ? tagArray_0_11 : _GEN_10; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_12 = 6'hc == CacheLineId ? tagArray_0_12 : _GEN_11; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_13 = 6'hd == CacheLineId ? tagArray_0_13 : _GEN_12; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_14 = 6'he == CacheLineId ? tagArray_0_14 : _GEN_13; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_15 = 6'hf == CacheLineId ? tagArray_0_15 : _GEN_14; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_16 = 6'h10 == CacheLineId ? tagArray_0_16 : _GEN_15; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_17 = 6'h11 == CacheLineId ? tagArray_0_17 : _GEN_16; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_18 = 6'h12 == CacheLineId ? tagArray_0_18 : _GEN_17; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_19 = 6'h13 == CacheLineId ? tagArray_0_19 : _GEN_18; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_20 = 6'h14 == CacheLineId ? tagArray_0_20 : _GEN_19; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_21 = 6'h15 == CacheLineId ? tagArray_0_21 : _GEN_20; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_22 = 6'h16 == CacheLineId ? tagArray_0_22 : _GEN_21; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_23 = 6'h17 == CacheLineId ? tagArray_0_23 : _GEN_22; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_24 = 6'h18 == CacheLineId ? tagArray_0_24 : _GEN_23; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_25 = 6'h19 == CacheLineId ? tagArray_0_25 : _GEN_24; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_26 = 6'h1a == CacheLineId ? tagArray_0_26 : _GEN_25; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_27 = 6'h1b == CacheLineId ? tagArray_0_27 : _GEN_26; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_28 = 6'h1c == CacheLineId ? tagArray_0_28 : _GEN_27; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_29 = 6'h1d == CacheLineId ? tagArray_0_29 : _GEN_28; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_30 = 6'h1e == CacheLineId ? tagArray_0_30 : _GEN_29; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_31 = 6'h1f == CacheLineId ? tagArray_0_31 : _GEN_30; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_32 = 6'h20 == CacheLineId ? tagArray_0_32 : _GEN_31; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_33 = 6'h21 == CacheLineId ? tagArray_0_33 : _GEN_32; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_34 = 6'h22 == CacheLineId ? tagArray_0_34 : _GEN_33; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_35 = 6'h23 == CacheLineId ? tagArray_0_35 : _GEN_34; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_36 = 6'h24 == CacheLineId ? tagArray_0_36 : _GEN_35; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_37 = 6'h25 == CacheLineId ? tagArray_0_37 : _GEN_36; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_38 = 6'h26 == CacheLineId ? tagArray_0_38 : _GEN_37; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_39 = 6'h27 == CacheLineId ? tagArray_0_39 : _GEN_38; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_40 = 6'h28 == CacheLineId ? tagArray_0_40 : _GEN_39; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_41 = 6'h29 == CacheLineId ? tagArray_0_41 : _GEN_40; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_42 = 6'h2a == CacheLineId ? tagArray_0_42 : _GEN_41; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_43 = 6'h2b == CacheLineId ? tagArray_0_43 : _GEN_42; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_44 = 6'h2c == CacheLineId ? tagArray_0_44 : _GEN_43; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_45 = 6'h2d == CacheLineId ? tagArray_0_45 : _GEN_44; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_46 = 6'h2e == CacheLineId ? tagArray_0_46 : _GEN_45; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_47 = 6'h2f == CacheLineId ? tagArray_0_47 : _GEN_46; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_48 = 6'h30 == CacheLineId ? tagArray_0_48 : _GEN_47; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_49 = 6'h31 == CacheLineId ? tagArray_0_49 : _GEN_48; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_50 = 6'h32 == CacheLineId ? tagArray_0_50 : _GEN_49; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_51 = 6'h33 == CacheLineId ? tagArray_0_51 : _GEN_50; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_52 = 6'h34 == CacheLineId ? tagArray_0_52 : _GEN_51; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_53 = 6'h35 == CacheLineId ? tagArray_0_53 : _GEN_52; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_54 = 6'h36 == CacheLineId ? tagArray_0_54 : _GEN_53; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_55 = 6'h37 == CacheLineId ? tagArray_0_55 : _GEN_54; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_56 = 6'h38 == CacheLineId ? tagArray_0_56 : _GEN_55; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_57 = 6'h39 == CacheLineId ? tagArray_0_57 : _GEN_56; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_58 = 6'h3a == CacheLineId ? tagArray_0_58 : _GEN_57; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_59 = 6'h3b == CacheLineId ? tagArray_0_59 : _GEN_58; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_60 = 6'h3c == CacheLineId ? tagArray_0_60 : _GEN_59; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_61 = 6'h3d == CacheLineId ? tagArray_0_61 : _GEN_60; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_62 = 6'h3e == CacheLineId ? tagArray_0_62 : _GEN_61; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_63 = 6'h3f == CacheLineId ? tagArray_0_63 : _GEN_62; // @[cache.scala 36:{14,14}]
  wire  _GEN_65 = 6'h1 == CacheLineId ? validArray_0_1 : validArray_0_0; // @[cache.scala 36:{44,44}]
  wire  _GEN_66 = 6'h2 == CacheLineId ? validArray_0_2 : _GEN_65; // @[cache.scala 36:{44,44}]
  wire  _GEN_67 = 6'h3 == CacheLineId ? validArray_0_3 : _GEN_66; // @[cache.scala 36:{44,44}]
  wire  _GEN_68 = 6'h4 == CacheLineId ? validArray_0_4 : _GEN_67; // @[cache.scala 36:{44,44}]
  wire  _GEN_69 = 6'h5 == CacheLineId ? validArray_0_5 : _GEN_68; // @[cache.scala 36:{44,44}]
  wire  _GEN_70 = 6'h6 == CacheLineId ? validArray_0_6 : _GEN_69; // @[cache.scala 36:{44,44}]
  wire  _GEN_71 = 6'h7 == CacheLineId ? validArray_0_7 : _GEN_70; // @[cache.scala 36:{44,44}]
  wire  _GEN_72 = 6'h8 == CacheLineId ? validArray_0_8 : _GEN_71; // @[cache.scala 36:{44,44}]
  wire  _GEN_73 = 6'h9 == CacheLineId ? validArray_0_9 : _GEN_72; // @[cache.scala 36:{44,44}]
  wire  _GEN_74 = 6'ha == CacheLineId ? validArray_0_10 : _GEN_73; // @[cache.scala 36:{44,44}]
  wire  _GEN_75 = 6'hb == CacheLineId ? validArray_0_11 : _GEN_74; // @[cache.scala 36:{44,44}]
  wire  _GEN_76 = 6'hc == CacheLineId ? validArray_0_12 : _GEN_75; // @[cache.scala 36:{44,44}]
  wire  _GEN_77 = 6'hd == CacheLineId ? validArray_0_13 : _GEN_76; // @[cache.scala 36:{44,44}]
  wire  _GEN_78 = 6'he == CacheLineId ? validArray_0_14 : _GEN_77; // @[cache.scala 36:{44,44}]
  wire  _GEN_79 = 6'hf == CacheLineId ? validArray_0_15 : _GEN_78; // @[cache.scala 36:{44,44}]
  wire  _GEN_80 = 6'h10 == CacheLineId ? validArray_0_16 : _GEN_79; // @[cache.scala 36:{44,44}]
  wire  _GEN_81 = 6'h11 == CacheLineId ? validArray_0_17 : _GEN_80; // @[cache.scala 36:{44,44}]
  wire  _GEN_82 = 6'h12 == CacheLineId ? validArray_0_18 : _GEN_81; // @[cache.scala 36:{44,44}]
  wire  _GEN_83 = 6'h13 == CacheLineId ? validArray_0_19 : _GEN_82; // @[cache.scala 36:{44,44}]
  wire  _GEN_84 = 6'h14 == CacheLineId ? validArray_0_20 : _GEN_83; // @[cache.scala 36:{44,44}]
  wire  _GEN_85 = 6'h15 == CacheLineId ? validArray_0_21 : _GEN_84; // @[cache.scala 36:{44,44}]
  wire  _GEN_86 = 6'h16 == CacheLineId ? validArray_0_22 : _GEN_85; // @[cache.scala 36:{44,44}]
  wire  _GEN_87 = 6'h17 == CacheLineId ? validArray_0_23 : _GEN_86; // @[cache.scala 36:{44,44}]
  wire  _GEN_88 = 6'h18 == CacheLineId ? validArray_0_24 : _GEN_87; // @[cache.scala 36:{44,44}]
  wire  _GEN_89 = 6'h19 == CacheLineId ? validArray_0_25 : _GEN_88; // @[cache.scala 36:{44,44}]
  wire  _GEN_90 = 6'h1a == CacheLineId ? validArray_0_26 : _GEN_89; // @[cache.scala 36:{44,44}]
  wire  _GEN_91 = 6'h1b == CacheLineId ? validArray_0_27 : _GEN_90; // @[cache.scala 36:{44,44}]
  wire  _GEN_92 = 6'h1c == CacheLineId ? validArray_0_28 : _GEN_91; // @[cache.scala 36:{44,44}]
  wire  _GEN_93 = 6'h1d == CacheLineId ? validArray_0_29 : _GEN_92; // @[cache.scala 36:{44,44}]
  wire  _GEN_94 = 6'h1e == CacheLineId ? validArray_0_30 : _GEN_93; // @[cache.scala 36:{44,44}]
  wire  _GEN_95 = 6'h1f == CacheLineId ? validArray_0_31 : _GEN_94; // @[cache.scala 36:{44,44}]
  wire  _GEN_96 = 6'h20 == CacheLineId ? validArray_0_32 : _GEN_95; // @[cache.scala 36:{44,44}]
  wire  _GEN_97 = 6'h21 == CacheLineId ? validArray_0_33 : _GEN_96; // @[cache.scala 36:{44,44}]
  wire  _GEN_98 = 6'h22 == CacheLineId ? validArray_0_34 : _GEN_97; // @[cache.scala 36:{44,44}]
  wire  _GEN_99 = 6'h23 == CacheLineId ? validArray_0_35 : _GEN_98; // @[cache.scala 36:{44,44}]
  wire  _GEN_100 = 6'h24 == CacheLineId ? validArray_0_36 : _GEN_99; // @[cache.scala 36:{44,44}]
  wire  _GEN_101 = 6'h25 == CacheLineId ? validArray_0_37 : _GEN_100; // @[cache.scala 36:{44,44}]
  wire  _GEN_102 = 6'h26 == CacheLineId ? validArray_0_38 : _GEN_101; // @[cache.scala 36:{44,44}]
  wire  _GEN_103 = 6'h27 == CacheLineId ? validArray_0_39 : _GEN_102; // @[cache.scala 36:{44,44}]
  wire  _GEN_104 = 6'h28 == CacheLineId ? validArray_0_40 : _GEN_103; // @[cache.scala 36:{44,44}]
  wire  _GEN_105 = 6'h29 == CacheLineId ? validArray_0_41 : _GEN_104; // @[cache.scala 36:{44,44}]
  wire  _GEN_106 = 6'h2a == CacheLineId ? validArray_0_42 : _GEN_105; // @[cache.scala 36:{44,44}]
  wire  _GEN_107 = 6'h2b == CacheLineId ? validArray_0_43 : _GEN_106; // @[cache.scala 36:{44,44}]
  wire  _GEN_108 = 6'h2c == CacheLineId ? validArray_0_44 : _GEN_107; // @[cache.scala 36:{44,44}]
  wire  _GEN_109 = 6'h2d == CacheLineId ? validArray_0_45 : _GEN_108; // @[cache.scala 36:{44,44}]
  wire  _GEN_110 = 6'h2e == CacheLineId ? validArray_0_46 : _GEN_109; // @[cache.scala 36:{44,44}]
  wire  _GEN_111 = 6'h2f == CacheLineId ? validArray_0_47 : _GEN_110; // @[cache.scala 36:{44,44}]
  wire  _GEN_112 = 6'h30 == CacheLineId ? validArray_0_48 : _GEN_111; // @[cache.scala 36:{44,44}]
  wire  _GEN_113 = 6'h31 == CacheLineId ? validArray_0_49 : _GEN_112; // @[cache.scala 36:{44,44}]
  wire  _GEN_114 = 6'h32 == CacheLineId ? validArray_0_50 : _GEN_113; // @[cache.scala 36:{44,44}]
  wire  _GEN_115 = 6'h33 == CacheLineId ? validArray_0_51 : _GEN_114; // @[cache.scala 36:{44,44}]
  wire  _GEN_116 = 6'h34 == CacheLineId ? validArray_0_52 : _GEN_115; // @[cache.scala 36:{44,44}]
  wire  _GEN_117 = 6'h35 == CacheLineId ? validArray_0_53 : _GEN_116; // @[cache.scala 36:{44,44}]
  wire  _GEN_118 = 6'h36 == CacheLineId ? validArray_0_54 : _GEN_117; // @[cache.scala 36:{44,44}]
  wire  _GEN_119 = 6'h37 == CacheLineId ? validArray_0_55 : _GEN_118; // @[cache.scala 36:{44,44}]
  wire  _GEN_120 = 6'h38 == CacheLineId ? validArray_0_56 : _GEN_119; // @[cache.scala 36:{44,44}]
  wire  _GEN_121 = 6'h39 == CacheLineId ? validArray_0_57 : _GEN_120; // @[cache.scala 36:{44,44}]
  wire  _GEN_122 = 6'h3a == CacheLineId ? validArray_0_58 : _GEN_121; // @[cache.scala 36:{44,44}]
  wire  _GEN_123 = 6'h3b == CacheLineId ? validArray_0_59 : _GEN_122; // @[cache.scala 36:{44,44}]
  wire  _GEN_124 = 6'h3c == CacheLineId ? validArray_0_60 : _GEN_123; // @[cache.scala 36:{44,44}]
  wire  _GEN_125 = 6'h3d == CacheLineId ? validArray_0_61 : _GEN_124; // @[cache.scala 36:{44,44}]
  wire  _GEN_126 = 6'h3e == CacheLineId ? validArray_0_62 : _GEN_125; // @[cache.scala 36:{44,44}]
  wire  _GEN_127 = 6'h3f == CacheLineId ? validArray_0_63 : _GEN_126; // @[cache.scala 36:{44,44}]
  wire  hitArray_0 = tag == _GEN_63 & _GEN_127; // @[cache.scala 36:44]
  wire [19:0] _GEN_129 = 6'h1 == CacheLineId ? tagArray_1_1 : tagArray_1_0; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_130 = 6'h2 == CacheLineId ? tagArray_1_2 : _GEN_129; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_131 = 6'h3 == CacheLineId ? tagArray_1_3 : _GEN_130; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_132 = 6'h4 == CacheLineId ? tagArray_1_4 : _GEN_131; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_133 = 6'h5 == CacheLineId ? tagArray_1_5 : _GEN_132; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_134 = 6'h6 == CacheLineId ? tagArray_1_6 : _GEN_133; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_135 = 6'h7 == CacheLineId ? tagArray_1_7 : _GEN_134; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_136 = 6'h8 == CacheLineId ? tagArray_1_8 : _GEN_135; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_137 = 6'h9 == CacheLineId ? tagArray_1_9 : _GEN_136; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_138 = 6'ha == CacheLineId ? tagArray_1_10 : _GEN_137; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_139 = 6'hb == CacheLineId ? tagArray_1_11 : _GEN_138; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_140 = 6'hc == CacheLineId ? tagArray_1_12 : _GEN_139; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_141 = 6'hd == CacheLineId ? tagArray_1_13 : _GEN_140; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_142 = 6'he == CacheLineId ? tagArray_1_14 : _GEN_141; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_143 = 6'hf == CacheLineId ? tagArray_1_15 : _GEN_142; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_144 = 6'h10 == CacheLineId ? tagArray_1_16 : _GEN_143; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_145 = 6'h11 == CacheLineId ? tagArray_1_17 : _GEN_144; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_146 = 6'h12 == CacheLineId ? tagArray_1_18 : _GEN_145; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_147 = 6'h13 == CacheLineId ? tagArray_1_19 : _GEN_146; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_148 = 6'h14 == CacheLineId ? tagArray_1_20 : _GEN_147; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_149 = 6'h15 == CacheLineId ? tagArray_1_21 : _GEN_148; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_150 = 6'h16 == CacheLineId ? tagArray_1_22 : _GEN_149; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_151 = 6'h17 == CacheLineId ? tagArray_1_23 : _GEN_150; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_152 = 6'h18 == CacheLineId ? tagArray_1_24 : _GEN_151; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_153 = 6'h19 == CacheLineId ? tagArray_1_25 : _GEN_152; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_154 = 6'h1a == CacheLineId ? tagArray_1_26 : _GEN_153; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_155 = 6'h1b == CacheLineId ? tagArray_1_27 : _GEN_154; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_156 = 6'h1c == CacheLineId ? tagArray_1_28 : _GEN_155; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_157 = 6'h1d == CacheLineId ? tagArray_1_29 : _GEN_156; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_158 = 6'h1e == CacheLineId ? tagArray_1_30 : _GEN_157; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_159 = 6'h1f == CacheLineId ? tagArray_1_31 : _GEN_158; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_160 = 6'h20 == CacheLineId ? tagArray_1_32 : _GEN_159; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_161 = 6'h21 == CacheLineId ? tagArray_1_33 : _GEN_160; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_162 = 6'h22 == CacheLineId ? tagArray_1_34 : _GEN_161; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_163 = 6'h23 == CacheLineId ? tagArray_1_35 : _GEN_162; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_164 = 6'h24 == CacheLineId ? tagArray_1_36 : _GEN_163; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_165 = 6'h25 == CacheLineId ? tagArray_1_37 : _GEN_164; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_166 = 6'h26 == CacheLineId ? tagArray_1_38 : _GEN_165; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_167 = 6'h27 == CacheLineId ? tagArray_1_39 : _GEN_166; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_168 = 6'h28 == CacheLineId ? tagArray_1_40 : _GEN_167; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_169 = 6'h29 == CacheLineId ? tagArray_1_41 : _GEN_168; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_170 = 6'h2a == CacheLineId ? tagArray_1_42 : _GEN_169; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_171 = 6'h2b == CacheLineId ? tagArray_1_43 : _GEN_170; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_172 = 6'h2c == CacheLineId ? tagArray_1_44 : _GEN_171; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_173 = 6'h2d == CacheLineId ? tagArray_1_45 : _GEN_172; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_174 = 6'h2e == CacheLineId ? tagArray_1_46 : _GEN_173; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_175 = 6'h2f == CacheLineId ? tagArray_1_47 : _GEN_174; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_176 = 6'h30 == CacheLineId ? tagArray_1_48 : _GEN_175; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_177 = 6'h31 == CacheLineId ? tagArray_1_49 : _GEN_176; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_178 = 6'h32 == CacheLineId ? tagArray_1_50 : _GEN_177; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_179 = 6'h33 == CacheLineId ? tagArray_1_51 : _GEN_178; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_180 = 6'h34 == CacheLineId ? tagArray_1_52 : _GEN_179; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_181 = 6'h35 == CacheLineId ? tagArray_1_53 : _GEN_180; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_182 = 6'h36 == CacheLineId ? tagArray_1_54 : _GEN_181; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_183 = 6'h37 == CacheLineId ? tagArray_1_55 : _GEN_182; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_184 = 6'h38 == CacheLineId ? tagArray_1_56 : _GEN_183; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_185 = 6'h39 == CacheLineId ? tagArray_1_57 : _GEN_184; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_186 = 6'h3a == CacheLineId ? tagArray_1_58 : _GEN_185; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_187 = 6'h3b == CacheLineId ? tagArray_1_59 : _GEN_186; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_188 = 6'h3c == CacheLineId ? tagArray_1_60 : _GEN_187; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_189 = 6'h3d == CacheLineId ? tagArray_1_61 : _GEN_188; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_190 = 6'h3e == CacheLineId ? tagArray_1_62 : _GEN_189; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_191 = 6'h3f == CacheLineId ? tagArray_1_63 : _GEN_190; // @[cache.scala 36:{14,14}]
  wire  _GEN_193 = 6'h1 == CacheLineId ? validArray_1_1 : validArray_1_0; // @[cache.scala 36:{44,44}]
  wire  _GEN_194 = 6'h2 == CacheLineId ? validArray_1_2 : _GEN_193; // @[cache.scala 36:{44,44}]
  wire  _GEN_195 = 6'h3 == CacheLineId ? validArray_1_3 : _GEN_194; // @[cache.scala 36:{44,44}]
  wire  _GEN_196 = 6'h4 == CacheLineId ? validArray_1_4 : _GEN_195; // @[cache.scala 36:{44,44}]
  wire  _GEN_197 = 6'h5 == CacheLineId ? validArray_1_5 : _GEN_196; // @[cache.scala 36:{44,44}]
  wire  _GEN_198 = 6'h6 == CacheLineId ? validArray_1_6 : _GEN_197; // @[cache.scala 36:{44,44}]
  wire  _GEN_199 = 6'h7 == CacheLineId ? validArray_1_7 : _GEN_198; // @[cache.scala 36:{44,44}]
  wire  _GEN_200 = 6'h8 == CacheLineId ? validArray_1_8 : _GEN_199; // @[cache.scala 36:{44,44}]
  wire  _GEN_201 = 6'h9 == CacheLineId ? validArray_1_9 : _GEN_200; // @[cache.scala 36:{44,44}]
  wire  _GEN_202 = 6'ha == CacheLineId ? validArray_1_10 : _GEN_201; // @[cache.scala 36:{44,44}]
  wire  _GEN_203 = 6'hb == CacheLineId ? validArray_1_11 : _GEN_202; // @[cache.scala 36:{44,44}]
  wire  _GEN_204 = 6'hc == CacheLineId ? validArray_1_12 : _GEN_203; // @[cache.scala 36:{44,44}]
  wire  _GEN_205 = 6'hd == CacheLineId ? validArray_1_13 : _GEN_204; // @[cache.scala 36:{44,44}]
  wire  _GEN_206 = 6'he == CacheLineId ? validArray_1_14 : _GEN_205; // @[cache.scala 36:{44,44}]
  wire  _GEN_207 = 6'hf == CacheLineId ? validArray_1_15 : _GEN_206; // @[cache.scala 36:{44,44}]
  wire  _GEN_208 = 6'h10 == CacheLineId ? validArray_1_16 : _GEN_207; // @[cache.scala 36:{44,44}]
  wire  _GEN_209 = 6'h11 == CacheLineId ? validArray_1_17 : _GEN_208; // @[cache.scala 36:{44,44}]
  wire  _GEN_210 = 6'h12 == CacheLineId ? validArray_1_18 : _GEN_209; // @[cache.scala 36:{44,44}]
  wire  _GEN_211 = 6'h13 == CacheLineId ? validArray_1_19 : _GEN_210; // @[cache.scala 36:{44,44}]
  wire  _GEN_212 = 6'h14 == CacheLineId ? validArray_1_20 : _GEN_211; // @[cache.scala 36:{44,44}]
  wire  _GEN_213 = 6'h15 == CacheLineId ? validArray_1_21 : _GEN_212; // @[cache.scala 36:{44,44}]
  wire  _GEN_214 = 6'h16 == CacheLineId ? validArray_1_22 : _GEN_213; // @[cache.scala 36:{44,44}]
  wire  _GEN_215 = 6'h17 == CacheLineId ? validArray_1_23 : _GEN_214; // @[cache.scala 36:{44,44}]
  wire  _GEN_216 = 6'h18 == CacheLineId ? validArray_1_24 : _GEN_215; // @[cache.scala 36:{44,44}]
  wire  _GEN_217 = 6'h19 == CacheLineId ? validArray_1_25 : _GEN_216; // @[cache.scala 36:{44,44}]
  wire  _GEN_218 = 6'h1a == CacheLineId ? validArray_1_26 : _GEN_217; // @[cache.scala 36:{44,44}]
  wire  _GEN_219 = 6'h1b == CacheLineId ? validArray_1_27 : _GEN_218; // @[cache.scala 36:{44,44}]
  wire  _GEN_220 = 6'h1c == CacheLineId ? validArray_1_28 : _GEN_219; // @[cache.scala 36:{44,44}]
  wire  _GEN_221 = 6'h1d == CacheLineId ? validArray_1_29 : _GEN_220; // @[cache.scala 36:{44,44}]
  wire  _GEN_222 = 6'h1e == CacheLineId ? validArray_1_30 : _GEN_221; // @[cache.scala 36:{44,44}]
  wire  _GEN_223 = 6'h1f == CacheLineId ? validArray_1_31 : _GEN_222; // @[cache.scala 36:{44,44}]
  wire  _GEN_224 = 6'h20 == CacheLineId ? validArray_1_32 : _GEN_223; // @[cache.scala 36:{44,44}]
  wire  _GEN_225 = 6'h21 == CacheLineId ? validArray_1_33 : _GEN_224; // @[cache.scala 36:{44,44}]
  wire  _GEN_226 = 6'h22 == CacheLineId ? validArray_1_34 : _GEN_225; // @[cache.scala 36:{44,44}]
  wire  _GEN_227 = 6'h23 == CacheLineId ? validArray_1_35 : _GEN_226; // @[cache.scala 36:{44,44}]
  wire  _GEN_228 = 6'h24 == CacheLineId ? validArray_1_36 : _GEN_227; // @[cache.scala 36:{44,44}]
  wire  _GEN_229 = 6'h25 == CacheLineId ? validArray_1_37 : _GEN_228; // @[cache.scala 36:{44,44}]
  wire  _GEN_230 = 6'h26 == CacheLineId ? validArray_1_38 : _GEN_229; // @[cache.scala 36:{44,44}]
  wire  _GEN_231 = 6'h27 == CacheLineId ? validArray_1_39 : _GEN_230; // @[cache.scala 36:{44,44}]
  wire  _GEN_232 = 6'h28 == CacheLineId ? validArray_1_40 : _GEN_231; // @[cache.scala 36:{44,44}]
  wire  _GEN_233 = 6'h29 == CacheLineId ? validArray_1_41 : _GEN_232; // @[cache.scala 36:{44,44}]
  wire  _GEN_234 = 6'h2a == CacheLineId ? validArray_1_42 : _GEN_233; // @[cache.scala 36:{44,44}]
  wire  _GEN_235 = 6'h2b == CacheLineId ? validArray_1_43 : _GEN_234; // @[cache.scala 36:{44,44}]
  wire  _GEN_236 = 6'h2c == CacheLineId ? validArray_1_44 : _GEN_235; // @[cache.scala 36:{44,44}]
  wire  _GEN_237 = 6'h2d == CacheLineId ? validArray_1_45 : _GEN_236; // @[cache.scala 36:{44,44}]
  wire  _GEN_238 = 6'h2e == CacheLineId ? validArray_1_46 : _GEN_237; // @[cache.scala 36:{44,44}]
  wire  _GEN_239 = 6'h2f == CacheLineId ? validArray_1_47 : _GEN_238; // @[cache.scala 36:{44,44}]
  wire  _GEN_240 = 6'h30 == CacheLineId ? validArray_1_48 : _GEN_239; // @[cache.scala 36:{44,44}]
  wire  _GEN_241 = 6'h31 == CacheLineId ? validArray_1_49 : _GEN_240; // @[cache.scala 36:{44,44}]
  wire  _GEN_242 = 6'h32 == CacheLineId ? validArray_1_50 : _GEN_241; // @[cache.scala 36:{44,44}]
  wire  _GEN_243 = 6'h33 == CacheLineId ? validArray_1_51 : _GEN_242; // @[cache.scala 36:{44,44}]
  wire  _GEN_244 = 6'h34 == CacheLineId ? validArray_1_52 : _GEN_243; // @[cache.scala 36:{44,44}]
  wire  _GEN_245 = 6'h35 == CacheLineId ? validArray_1_53 : _GEN_244; // @[cache.scala 36:{44,44}]
  wire  _GEN_246 = 6'h36 == CacheLineId ? validArray_1_54 : _GEN_245; // @[cache.scala 36:{44,44}]
  wire  _GEN_247 = 6'h37 == CacheLineId ? validArray_1_55 : _GEN_246; // @[cache.scala 36:{44,44}]
  wire  _GEN_248 = 6'h38 == CacheLineId ? validArray_1_56 : _GEN_247; // @[cache.scala 36:{44,44}]
  wire  _GEN_249 = 6'h39 == CacheLineId ? validArray_1_57 : _GEN_248; // @[cache.scala 36:{44,44}]
  wire  _GEN_250 = 6'h3a == CacheLineId ? validArray_1_58 : _GEN_249; // @[cache.scala 36:{44,44}]
  wire  _GEN_251 = 6'h3b == CacheLineId ? validArray_1_59 : _GEN_250; // @[cache.scala 36:{44,44}]
  wire  _GEN_252 = 6'h3c == CacheLineId ? validArray_1_60 : _GEN_251; // @[cache.scala 36:{44,44}]
  wire  _GEN_253 = 6'h3d == CacheLineId ? validArray_1_61 : _GEN_252; // @[cache.scala 36:{44,44}]
  wire  _GEN_254 = 6'h3e == CacheLineId ? validArray_1_62 : _GEN_253; // @[cache.scala 36:{44,44}]
  wire  _GEN_255 = 6'h3f == CacheLineId ? validArray_1_63 : _GEN_254; // @[cache.scala 36:{44,44}]
  wire  hitArray_1 = tag == _GEN_191 & _GEN_255; // @[cache.scala 36:44]
  wire [19:0] _GEN_257 = 6'h1 == CacheLineId ? tagArray_2_1 : tagArray_2_0; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_258 = 6'h2 == CacheLineId ? tagArray_2_2 : _GEN_257; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_259 = 6'h3 == CacheLineId ? tagArray_2_3 : _GEN_258; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_260 = 6'h4 == CacheLineId ? tagArray_2_4 : _GEN_259; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_261 = 6'h5 == CacheLineId ? tagArray_2_5 : _GEN_260; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_262 = 6'h6 == CacheLineId ? tagArray_2_6 : _GEN_261; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_263 = 6'h7 == CacheLineId ? tagArray_2_7 : _GEN_262; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_264 = 6'h8 == CacheLineId ? tagArray_2_8 : _GEN_263; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_265 = 6'h9 == CacheLineId ? tagArray_2_9 : _GEN_264; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_266 = 6'ha == CacheLineId ? tagArray_2_10 : _GEN_265; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_267 = 6'hb == CacheLineId ? tagArray_2_11 : _GEN_266; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_268 = 6'hc == CacheLineId ? tagArray_2_12 : _GEN_267; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_269 = 6'hd == CacheLineId ? tagArray_2_13 : _GEN_268; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_270 = 6'he == CacheLineId ? tagArray_2_14 : _GEN_269; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_271 = 6'hf == CacheLineId ? tagArray_2_15 : _GEN_270; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_272 = 6'h10 == CacheLineId ? tagArray_2_16 : _GEN_271; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_273 = 6'h11 == CacheLineId ? tagArray_2_17 : _GEN_272; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_274 = 6'h12 == CacheLineId ? tagArray_2_18 : _GEN_273; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_275 = 6'h13 == CacheLineId ? tagArray_2_19 : _GEN_274; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_276 = 6'h14 == CacheLineId ? tagArray_2_20 : _GEN_275; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_277 = 6'h15 == CacheLineId ? tagArray_2_21 : _GEN_276; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_278 = 6'h16 == CacheLineId ? tagArray_2_22 : _GEN_277; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_279 = 6'h17 == CacheLineId ? tagArray_2_23 : _GEN_278; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_280 = 6'h18 == CacheLineId ? tagArray_2_24 : _GEN_279; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_281 = 6'h19 == CacheLineId ? tagArray_2_25 : _GEN_280; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_282 = 6'h1a == CacheLineId ? tagArray_2_26 : _GEN_281; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_283 = 6'h1b == CacheLineId ? tagArray_2_27 : _GEN_282; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_284 = 6'h1c == CacheLineId ? tagArray_2_28 : _GEN_283; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_285 = 6'h1d == CacheLineId ? tagArray_2_29 : _GEN_284; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_286 = 6'h1e == CacheLineId ? tagArray_2_30 : _GEN_285; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_287 = 6'h1f == CacheLineId ? tagArray_2_31 : _GEN_286; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_288 = 6'h20 == CacheLineId ? tagArray_2_32 : _GEN_287; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_289 = 6'h21 == CacheLineId ? tagArray_2_33 : _GEN_288; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_290 = 6'h22 == CacheLineId ? tagArray_2_34 : _GEN_289; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_291 = 6'h23 == CacheLineId ? tagArray_2_35 : _GEN_290; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_292 = 6'h24 == CacheLineId ? tagArray_2_36 : _GEN_291; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_293 = 6'h25 == CacheLineId ? tagArray_2_37 : _GEN_292; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_294 = 6'h26 == CacheLineId ? tagArray_2_38 : _GEN_293; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_295 = 6'h27 == CacheLineId ? tagArray_2_39 : _GEN_294; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_296 = 6'h28 == CacheLineId ? tagArray_2_40 : _GEN_295; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_297 = 6'h29 == CacheLineId ? tagArray_2_41 : _GEN_296; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_298 = 6'h2a == CacheLineId ? tagArray_2_42 : _GEN_297; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_299 = 6'h2b == CacheLineId ? tagArray_2_43 : _GEN_298; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_300 = 6'h2c == CacheLineId ? tagArray_2_44 : _GEN_299; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_301 = 6'h2d == CacheLineId ? tagArray_2_45 : _GEN_300; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_302 = 6'h2e == CacheLineId ? tagArray_2_46 : _GEN_301; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_303 = 6'h2f == CacheLineId ? tagArray_2_47 : _GEN_302; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_304 = 6'h30 == CacheLineId ? tagArray_2_48 : _GEN_303; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_305 = 6'h31 == CacheLineId ? tagArray_2_49 : _GEN_304; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_306 = 6'h32 == CacheLineId ? tagArray_2_50 : _GEN_305; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_307 = 6'h33 == CacheLineId ? tagArray_2_51 : _GEN_306; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_308 = 6'h34 == CacheLineId ? tagArray_2_52 : _GEN_307; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_309 = 6'h35 == CacheLineId ? tagArray_2_53 : _GEN_308; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_310 = 6'h36 == CacheLineId ? tagArray_2_54 : _GEN_309; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_311 = 6'h37 == CacheLineId ? tagArray_2_55 : _GEN_310; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_312 = 6'h38 == CacheLineId ? tagArray_2_56 : _GEN_311; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_313 = 6'h39 == CacheLineId ? tagArray_2_57 : _GEN_312; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_314 = 6'h3a == CacheLineId ? tagArray_2_58 : _GEN_313; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_315 = 6'h3b == CacheLineId ? tagArray_2_59 : _GEN_314; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_316 = 6'h3c == CacheLineId ? tagArray_2_60 : _GEN_315; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_317 = 6'h3d == CacheLineId ? tagArray_2_61 : _GEN_316; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_318 = 6'h3e == CacheLineId ? tagArray_2_62 : _GEN_317; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_319 = 6'h3f == CacheLineId ? tagArray_2_63 : _GEN_318; // @[cache.scala 36:{14,14}]
  wire  _GEN_321 = 6'h1 == CacheLineId ? validArray_2_1 : validArray_2_0; // @[cache.scala 36:{44,44}]
  wire  _GEN_322 = 6'h2 == CacheLineId ? validArray_2_2 : _GEN_321; // @[cache.scala 36:{44,44}]
  wire  _GEN_323 = 6'h3 == CacheLineId ? validArray_2_3 : _GEN_322; // @[cache.scala 36:{44,44}]
  wire  _GEN_324 = 6'h4 == CacheLineId ? validArray_2_4 : _GEN_323; // @[cache.scala 36:{44,44}]
  wire  _GEN_325 = 6'h5 == CacheLineId ? validArray_2_5 : _GEN_324; // @[cache.scala 36:{44,44}]
  wire  _GEN_326 = 6'h6 == CacheLineId ? validArray_2_6 : _GEN_325; // @[cache.scala 36:{44,44}]
  wire  _GEN_327 = 6'h7 == CacheLineId ? validArray_2_7 : _GEN_326; // @[cache.scala 36:{44,44}]
  wire  _GEN_328 = 6'h8 == CacheLineId ? validArray_2_8 : _GEN_327; // @[cache.scala 36:{44,44}]
  wire  _GEN_329 = 6'h9 == CacheLineId ? validArray_2_9 : _GEN_328; // @[cache.scala 36:{44,44}]
  wire  _GEN_330 = 6'ha == CacheLineId ? validArray_2_10 : _GEN_329; // @[cache.scala 36:{44,44}]
  wire  _GEN_331 = 6'hb == CacheLineId ? validArray_2_11 : _GEN_330; // @[cache.scala 36:{44,44}]
  wire  _GEN_332 = 6'hc == CacheLineId ? validArray_2_12 : _GEN_331; // @[cache.scala 36:{44,44}]
  wire  _GEN_333 = 6'hd == CacheLineId ? validArray_2_13 : _GEN_332; // @[cache.scala 36:{44,44}]
  wire  _GEN_334 = 6'he == CacheLineId ? validArray_2_14 : _GEN_333; // @[cache.scala 36:{44,44}]
  wire  _GEN_335 = 6'hf == CacheLineId ? validArray_2_15 : _GEN_334; // @[cache.scala 36:{44,44}]
  wire  _GEN_336 = 6'h10 == CacheLineId ? validArray_2_16 : _GEN_335; // @[cache.scala 36:{44,44}]
  wire  _GEN_337 = 6'h11 == CacheLineId ? validArray_2_17 : _GEN_336; // @[cache.scala 36:{44,44}]
  wire  _GEN_338 = 6'h12 == CacheLineId ? validArray_2_18 : _GEN_337; // @[cache.scala 36:{44,44}]
  wire  _GEN_339 = 6'h13 == CacheLineId ? validArray_2_19 : _GEN_338; // @[cache.scala 36:{44,44}]
  wire  _GEN_340 = 6'h14 == CacheLineId ? validArray_2_20 : _GEN_339; // @[cache.scala 36:{44,44}]
  wire  _GEN_341 = 6'h15 == CacheLineId ? validArray_2_21 : _GEN_340; // @[cache.scala 36:{44,44}]
  wire  _GEN_342 = 6'h16 == CacheLineId ? validArray_2_22 : _GEN_341; // @[cache.scala 36:{44,44}]
  wire  _GEN_343 = 6'h17 == CacheLineId ? validArray_2_23 : _GEN_342; // @[cache.scala 36:{44,44}]
  wire  _GEN_344 = 6'h18 == CacheLineId ? validArray_2_24 : _GEN_343; // @[cache.scala 36:{44,44}]
  wire  _GEN_345 = 6'h19 == CacheLineId ? validArray_2_25 : _GEN_344; // @[cache.scala 36:{44,44}]
  wire  _GEN_346 = 6'h1a == CacheLineId ? validArray_2_26 : _GEN_345; // @[cache.scala 36:{44,44}]
  wire  _GEN_347 = 6'h1b == CacheLineId ? validArray_2_27 : _GEN_346; // @[cache.scala 36:{44,44}]
  wire  _GEN_348 = 6'h1c == CacheLineId ? validArray_2_28 : _GEN_347; // @[cache.scala 36:{44,44}]
  wire  _GEN_349 = 6'h1d == CacheLineId ? validArray_2_29 : _GEN_348; // @[cache.scala 36:{44,44}]
  wire  _GEN_350 = 6'h1e == CacheLineId ? validArray_2_30 : _GEN_349; // @[cache.scala 36:{44,44}]
  wire  _GEN_351 = 6'h1f == CacheLineId ? validArray_2_31 : _GEN_350; // @[cache.scala 36:{44,44}]
  wire  _GEN_352 = 6'h20 == CacheLineId ? validArray_2_32 : _GEN_351; // @[cache.scala 36:{44,44}]
  wire  _GEN_353 = 6'h21 == CacheLineId ? validArray_2_33 : _GEN_352; // @[cache.scala 36:{44,44}]
  wire  _GEN_354 = 6'h22 == CacheLineId ? validArray_2_34 : _GEN_353; // @[cache.scala 36:{44,44}]
  wire  _GEN_355 = 6'h23 == CacheLineId ? validArray_2_35 : _GEN_354; // @[cache.scala 36:{44,44}]
  wire  _GEN_356 = 6'h24 == CacheLineId ? validArray_2_36 : _GEN_355; // @[cache.scala 36:{44,44}]
  wire  _GEN_357 = 6'h25 == CacheLineId ? validArray_2_37 : _GEN_356; // @[cache.scala 36:{44,44}]
  wire  _GEN_358 = 6'h26 == CacheLineId ? validArray_2_38 : _GEN_357; // @[cache.scala 36:{44,44}]
  wire  _GEN_359 = 6'h27 == CacheLineId ? validArray_2_39 : _GEN_358; // @[cache.scala 36:{44,44}]
  wire  _GEN_360 = 6'h28 == CacheLineId ? validArray_2_40 : _GEN_359; // @[cache.scala 36:{44,44}]
  wire  _GEN_361 = 6'h29 == CacheLineId ? validArray_2_41 : _GEN_360; // @[cache.scala 36:{44,44}]
  wire  _GEN_362 = 6'h2a == CacheLineId ? validArray_2_42 : _GEN_361; // @[cache.scala 36:{44,44}]
  wire  _GEN_363 = 6'h2b == CacheLineId ? validArray_2_43 : _GEN_362; // @[cache.scala 36:{44,44}]
  wire  _GEN_364 = 6'h2c == CacheLineId ? validArray_2_44 : _GEN_363; // @[cache.scala 36:{44,44}]
  wire  _GEN_365 = 6'h2d == CacheLineId ? validArray_2_45 : _GEN_364; // @[cache.scala 36:{44,44}]
  wire  _GEN_366 = 6'h2e == CacheLineId ? validArray_2_46 : _GEN_365; // @[cache.scala 36:{44,44}]
  wire  _GEN_367 = 6'h2f == CacheLineId ? validArray_2_47 : _GEN_366; // @[cache.scala 36:{44,44}]
  wire  _GEN_368 = 6'h30 == CacheLineId ? validArray_2_48 : _GEN_367; // @[cache.scala 36:{44,44}]
  wire  _GEN_369 = 6'h31 == CacheLineId ? validArray_2_49 : _GEN_368; // @[cache.scala 36:{44,44}]
  wire  _GEN_370 = 6'h32 == CacheLineId ? validArray_2_50 : _GEN_369; // @[cache.scala 36:{44,44}]
  wire  _GEN_371 = 6'h33 == CacheLineId ? validArray_2_51 : _GEN_370; // @[cache.scala 36:{44,44}]
  wire  _GEN_372 = 6'h34 == CacheLineId ? validArray_2_52 : _GEN_371; // @[cache.scala 36:{44,44}]
  wire  _GEN_373 = 6'h35 == CacheLineId ? validArray_2_53 : _GEN_372; // @[cache.scala 36:{44,44}]
  wire  _GEN_374 = 6'h36 == CacheLineId ? validArray_2_54 : _GEN_373; // @[cache.scala 36:{44,44}]
  wire  _GEN_375 = 6'h37 == CacheLineId ? validArray_2_55 : _GEN_374; // @[cache.scala 36:{44,44}]
  wire  _GEN_376 = 6'h38 == CacheLineId ? validArray_2_56 : _GEN_375; // @[cache.scala 36:{44,44}]
  wire  _GEN_377 = 6'h39 == CacheLineId ? validArray_2_57 : _GEN_376; // @[cache.scala 36:{44,44}]
  wire  _GEN_378 = 6'h3a == CacheLineId ? validArray_2_58 : _GEN_377; // @[cache.scala 36:{44,44}]
  wire  _GEN_379 = 6'h3b == CacheLineId ? validArray_2_59 : _GEN_378; // @[cache.scala 36:{44,44}]
  wire  _GEN_380 = 6'h3c == CacheLineId ? validArray_2_60 : _GEN_379; // @[cache.scala 36:{44,44}]
  wire  _GEN_381 = 6'h3d == CacheLineId ? validArray_2_61 : _GEN_380; // @[cache.scala 36:{44,44}]
  wire  _GEN_382 = 6'h3e == CacheLineId ? validArray_2_62 : _GEN_381; // @[cache.scala 36:{44,44}]
  wire  _GEN_383 = 6'h3f == CacheLineId ? validArray_2_63 : _GEN_382; // @[cache.scala 36:{44,44}]
  wire  hitArray_2 = tag == _GEN_319 & _GEN_383; // @[cache.scala 36:44]
  wire [19:0] _GEN_385 = 6'h1 == CacheLineId ? tagArray_3_1 : tagArray_3_0; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_386 = 6'h2 == CacheLineId ? tagArray_3_2 : _GEN_385; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_387 = 6'h3 == CacheLineId ? tagArray_3_3 : _GEN_386; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_388 = 6'h4 == CacheLineId ? tagArray_3_4 : _GEN_387; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_389 = 6'h5 == CacheLineId ? tagArray_3_5 : _GEN_388; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_390 = 6'h6 == CacheLineId ? tagArray_3_6 : _GEN_389; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_391 = 6'h7 == CacheLineId ? tagArray_3_7 : _GEN_390; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_392 = 6'h8 == CacheLineId ? tagArray_3_8 : _GEN_391; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_393 = 6'h9 == CacheLineId ? tagArray_3_9 : _GEN_392; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_394 = 6'ha == CacheLineId ? tagArray_3_10 : _GEN_393; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_395 = 6'hb == CacheLineId ? tagArray_3_11 : _GEN_394; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_396 = 6'hc == CacheLineId ? tagArray_3_12 : _GEN_395; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_397 = 6'hd == CacheLineId ? tagArray_3_13 : _GEN_396; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_398 = 6'he == CacheLineId ? tagArray_3_14 : _GEN_397; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_399 = 6'hf == CacheLineId ? tagArray_3_15 : _GEN_398; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_400 = 6'h10 == CacheLineId ? tagArray_3_16 : _GEN_399; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_401 = 6'h11 == CacheLineId ? tagArray_3_17 : _GEN_400; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_402 = 6'h12 == CacheLineId ? tagArray_3_18 : _GEN_401; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_403 = 6'h13 == CacheLineId ? tagArray_3_19 : _GEN_402; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_404 = 6'h14 == CacheLineId ? tagArray_3_20 : _GEN_403; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_405 = 6'h15 == CacheLineId ? tagArray_3_21 : _GEN_404; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_406 = 6'h16 == CacheLineId ? tagArray_3_22 : _GEN_405; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_407 = 6'h17 == CacheLineId ? tagArray_3_23 : _GEN_406; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_408 = 6'h18 == CacheLineId ? tagArray_3_24 : _GEN_407; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_409 = 6'h19 == CacheLineId ? tagArray_3_25 : _GEN_408; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_410 = 6'h1a == CacheLineId ? tagArray_3_26 : _GEN_409; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_411 = 6'h1b == CacheLineId ? tagArray_3_27 : _GEN_410; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_412 = 6'h1c == CacheLineId ? tagArray_3_28 : _GEN_411; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_413 = 6'h1d == CacheLineId ? tagArray_3_29 : _GEN_412; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_414 = 6'h1e == CacheLineId ? tagArray_3_30 : _GEN_413; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_415 = 6'h1f == CacheLineId ? tagArray_3_31 : _GEN_414; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_416 = 6'h20 == CacheLineId ? tagArray_3_32 : _GEN_415; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_417 = 6'h21 == CacheLineId ? tagArray_3_33 : _GEN_416; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_418 = 6'h22 == CacheLineId ? tagArray_3_34 : _GEN_417; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_419 = 6'h23 == CacheLineId ? tagArray_3_35 : _GEN_418; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_420 = 6'h24 == CacheLineId ? tagArray_3_36 : _GEN_419; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_421 = 6'h25 == CacheLineId ? tagArray_3_37 : _GEN_420; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_422 = 6'h26 == CacheLineId ? tagArray_3_38 : _GEN_421; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_423 = 6'h27 == CacheLineId ? tagArray_3_39 : _GEN_422; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_424 = 6'h28 == CacheLineId ? tagArray_3_40 : _GEN_423; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_425 = 6'h29 == CacheLineId ? tagArray_3_41 : _GEN_424; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_426 = 6'h2a == CacheLineId ? tagArray_3_42 : _GEN_425; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_427 = 6'h2b == CacheLineId ? tagArray_3_43 : _GEN_426; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_428 = 6'h2c == CacheLineId ? tagArray_3_44 : _GEN_427; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_429 = 6'h2d == CacheLineId ? tagArray_3_45 : _GEN_428; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_430 = 6'h2e == CacheLineId ? tagArray_3_46 : _GEN_429; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_431 = 6'h2f == CacheLineId ? tagArray_3_47 : _GEN_430; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_432 = 6'h30 == CacheLineId ? tagArray_3_48 : _GEN_431; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_433 = 6'h31 == CacheLineId ? tagArray_3_49 : _GEN_432; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_434 = 6'h32 == CacheLineId ? tagArray_3_50 : _GEN_433; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_435 = 6'h33 == CacheLineId ? tagArray_3_51 : _GEN_434; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_436 = 6'h34 == CacheLineId ? tagArray_3_52 : _GEN_435; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_437 = 6'h35 == CacheLineId ? tagArray_3_53 : _GEN_436; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_438 = 6'h36 == CacheLineId ? tagArray_3_54 : _GEN_437; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_439 = 6'h37 == CacheLineId ? tagArray_3_55 : _GEN_438; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_440 = 6'h38 == CacheLineId ? tagArray_3_56 : _GEN_439; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_441 = 6'h39 == CacheLineId ? tagArray_3_57 : _GEN_440; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_442 = 6'h3a == CacheLineId ? tagArray_3_58 : _GEN_441; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_443 = 6'h3b == CacheLineId ? tagArray_3_59 : _GEN_442; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_444 = 6'h3c == CacheLineId ? tagArray_3_60 : _GEN_443; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_445 = 6'h3d == CacheLineId ? tagArray_3_61 : _GEN_444; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_446 = 6'h3e == CacheLineId ? tagArray_3_62 : _GEN_445; // @[cache.scala 36:{14,14}]
  wire [19:0] _GEN_447 = 6'h3f == CacheLineId ? tagArray_3_63 : _GEN_446; // @[cache.scala 36:{14,14}]
  wire  _GEN_449 = 6'h1 == CacheLineId ? validArray_3_1 : validArray_3_0; // @[cache.scala 36:{44,44}]
  wire  _GEN_450 = 6'h2 == CacheLineId ? validArray_3_2 : _GEN_449; // @[cache.scala 36:{44,44}]
  wire  _GEN_451 = 6'h3 == CacheLineId ? validArray_3_3 : _GEN_450; // @[cache.scala 36:{44,44}]
  wire  _GEN_452 = 6'h4 == CacheLineId ? validArray_3_4 : _GEN_451; // @[cache.scala 36:{44,44}]
  wire  _GEN_453 = 6'h5 == CacheLineId ? validArray_3_5 : _GEN_452; // @[cache.scala 36:{44,44}]
  wire  _GEN_454 = 6'h6 == CacheLineId ? validArray_3_6 : _GEN_453; // @[cache.scala 36:{44,44}]
  wire  _GEN_455 = 6'h7 == CacheLineId ? validArray_3_7 : _GEN_454; // @[cache.scala 36:{44,44}]
  wire  _GEN_456 = 6'h8 == CacheLineId ? validArray_3_8 : _GEN_455; // @[cache.scala 36:{44,44}]
  wire  _GEN_457 = 6'h9 == CacheLineId ? validArray_3_9 : _GEN_456; // @[cache.scala 36:{44,44}]
  wire  _GEN_458 = 6'ha == CacheLineId ? validArray_3_10 : _GEN_457; // @[cache.scala 36:{44,44}]
  wire  _GEN_459 = 6'hb == CacheLineId ? validArray_3_11 : _GEN_458; // @[cache.scala 36:{44,44}]
  wire  _GEN_460 = 6'hc == CacheLineId ? validArray_3_12 : _GEN_459; // @[cache.scala 36:{44,44}]
  wire  _GEN_461 = 6'hd == CacheLineId ? validArray_3_13 : _GEN_460; // @[cache.scala 36:{44,44}]
  wire  _GEN_462 = 6'he == CacheLineId ? validArray_3_14 : _GEN_461; // @[cache.scala 36:{44,44}]
  wire  _GEN_463 = 6'hf == CacheLineId ? validArray_3_15 : _GEN_462; // @[cache.scala 36:{44,44}]
  wire  _GEN_464 = 6'h10 == CacheLineId ? validArray_3_16 : _GEN_463; // @[cache.scala 36:{44,44}]
  wire  _GEN_465 = 6'h11 == CacheLineId ? validArray_3_17 : _GEN_464; // @[cache.scala 36:{44,44}]
  wire  _GEN_466 = 6'h12 == CacheLineId ? validArray_3_18 : _GEN_465; // @[cache.scala 36:{44,44}]
  wire  _GEN_467 = 6'h13 == CacheLineId ? validArray_3_19 : _GEN_466; // @[cache.scala 36:{44,44}]
  wire  _GEN_468 = 6'h14 == CacheLineId ? validArray_3_20 : _GEN_467; // @[cache.scala 36:{44,44}]
  wire  _GEN_469 = 6'h15 == CacheLineId ? validArray_3_21 : _GEN_468; // @[cache.scala 36:{44,44}]
  wire  _GEN_470 = 6'h16 == CacheLineId ? validArray_3_22 : _GEN_469; // @[cache.scala 36:{44,44}]
  wire  _GEN_471 = 6'h17 == CacheLineId ? validArray_3_23 : _GEN_470; // @[cache.scala 36:{44,44}]
  wire  _GEN_472 = 6'h18 == CacheLineId ? validArray_3_24 : _GEN_471; // @[cache.scala 36:{44,44}]
  wire  _GEN_473 = 6'h19 == CacheLineId ? validArray_3_25 : _GEN_472; // @[cache.scala 36:{44,44}]
  wire  _GEN_474 = 6'h1a == CacheLineId ? validArray_3_26 : _GEN_473; // @[cache.scala 36:{44,44}]
  wire  _GEN_475 = 6'h1b == CacheLineId ? validArray_3_27 : _GEN_474; // @[cache.scala 36:{44,44}]
  wire  _GEN_476 = 6'h1c == CacheLineId ? validArray_3_28 : _GEN_475; // @[cache.scala 36:{44,44}]
  wire  _GEN_477 = 6'h1d == CacheLineId ? validArray_3_29 : _GEN_476; // @[cache.scala 36:{44,44}]
  wire  _GEN_478 = 6'h1e == CacheLineId ? validArray_3_30 : _GEN_477; // @[cache.scala 36:{44,44}]
  wire  _GEN_479 = 6'h1f == CacheLineId ? validArray_3_31 : _GEN_478; // @[cache.scala 36:{44,44}]
  wire  _GEN_480 = 6'h20 == CacheLineId ? validArray_3_32 : _GEN_479; // @[cache.scala 36:{44,44}]
  wire  _GEN_481 = 6'h21 == CacheLineId ? validArray_3_33 : _GEN_480; // @[cache.scala 36:{44,44}]
  wire  _GEN_482 = 6'h22 == CacheLineId ? validArray_3_34 : _GEN_481; // @[cache.scala 36:{44,44}]
  wire  _GEN_483 = 6'h23 == CacheLineId ? validArray_3_35 : _GEN_482; // @[cache.scala 36:{44,44}]
  wire  _GEN_484 = 6'h24 == CacheLineId ? validArray_3_36 : _GEN_483; // @[cache.scala 36:{44,44}]
  wire  _GEN_485 = 6'h25 == CacheLineId ? validArray_3_37 : _GEN_484; // @[cache.scala 36:{44,44}]
  wire  _GEN_486 = 6'h26 == CacheLineId ? validArray_3_38 : _GEN_485; // @[cache.scala 36:{44,44}]
  wire  _GEN_487 = 6'h27 == CacheLineId ? validArray_3_39 : _GEN_486; // @[cache.scala 36:{44,44}]
  wire  _GEN_488 = 6'h28 == CacheLineId ? validArray_3_40 : _GEN_487; // @[cache.scala 36:{44,44}]
  wire  _GEN_489 = 6'h29 == CacheLineId ? validArray_3_41 : _GEN_488; // @[cache.scala 36:{44,44}]
  wire  _GEN_490 = 6'h2a == CacheLineId ? validArray_3_42 : _GEN_489; // @[cache.scala 36:{44,44}]
  wire  _GEN_491 = 6'h2b == CacheLineId ? validArray_3_43 : _GEN_490; // @[cache.scala 36:{44,44}]
  wire  _GEN_492 = 6'h2c == CacheLineId ? validArray_3_44 : _GEN_491; // @[cache.scala 36:{44,44}]
  wire  _GEN_493 = 6'h2d == CacheLineId ? validArray_3_45 : _GEN_492; // @[cache.scala 36:{44,44}]
  wire  _GEN_494 = 6'h2e == CacheLineId ? validArray_3_46 : _GEN_493; // @[cache.scala 36:{44,44}]
  wire  _GEN_495 = 6'h2f == CacheLineId ? validArray_3_47 : _GEN_494; // @[cache.scala 36:{44,44}]
  wire  _GEN_496 = 6'h30 == CacheLineId ? validArray_3_48 : _GEN_495; // @[cache.scala 36:{44,44}]
  wire  _GEN_497 = 6'h31 == CacheLineId ? validArray_3_49 : _GEN_496; // @[cache.scala 36:{44,44}]
  wire  _GEN_498 = 6'h32 == CacheLineId ? validArray_3_50 : _GEN_497; // @[cache.scala 36:{44,44}]
  wire  _GEN_499 = 6'h33 == CacheLineId ? validArray_3_51 : _GEN_498; // @[cache.scala 36:{44,44}]
  wire  _GEN_500 = 6'h34 == CacheLineId ? validArray_3_52 : _GEN_499; // @[cache.scala 36:{44,44}]
  wire  _GEN_501 = 6'h35 == CacheLineId ? validArray_3_53 : _GEN_500; // @[cache.scala 36:{44,44}]
  wire  _GEN_502 = 6'h36 == CacheLineId ? validArray_3_54 : _GEN_501; // @[cache.scala 36:{44,44}]
  wire  _GEN_503 = 6'h37 == CacheLineId ? validArray_3_55 : _GEN_502; // @[cache.scala 36:{44,44}]
  wire  _GEN_504 = 6'h38 == CacheLineId ? validArray_3_56 : _GEN_503; // @[cache.scala 36:{44,44}]
  wire  _GEN_505 = 6'h39 == CacheLineId ? validArray_3_57 : _GEN_504; // @[cache.scala 36:{44,44}]
  wire  _GEN_506 = 6'h3a == CacheLineId ? validArray_3_58 : _GEN_505; // @[cache.scala 36:{44,44}]
  wire  _GEN_507 = 6'h3b == CacheLineId ? validArray_3_59 : _GEN_506; // @[cache.scala 36:{44,44}]
  wire  _GEN_508 = 6'h3c == CacheLineId ? validArray_3_60 : _GEN_507; // @[cache.scala 36:{44,44}]
  wire  _GEN_509 = 6'h3d == CacheLineId ? validArray_3_61 : _GEN_508; // @[cache.scala 36:{44,44}]
  wire  _GEN_510 = 6'h3e == CacheLineId ? validArray_3_62 : _GEN_509; // @[cache.scala 36:{44,44}]
  wire  _GEN_511 = 6'h3f == CacheLineId ? validArray_3_63 : _GEN_510; // @[cache.scala 36:{44,44}]
  wire  hitArray_3 = tag == _GEN_447 & _GEN_511; // @[cache.scala 36:44]
  wire  hit = hitArray_0 | hitArray_1 | hitArray_2 | hitArray_3; // @[cache.scala 38:33]
  wire  _SetId_T_6 = _GEN_447 == tag; // @[Mux.scala 81:61]
  reg [3:0] off; // @[cache.scala 45:24]
  reg [2:0] state_cache; // @[cache.scala 48:30]
  wire  _T_1 = from_IFU_ready & from_IFU_valid; // @[Decoupled.scala 51:35]
  wire  _T_3 = 3'h2 == state_cache; // @[cache.scala 49:26]
  wire  _state_cache_T_1 = to_sram_ar_ready & to_sram_ar_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_cache_T_2 = _state_cache_T_1 ? 3'h3 : 3'h2; // @[cache.scala 62:31]
  wire [2:0] _state_cache_T_3 = to_sram_r_bits_last ? 3'h4 : 3'h3; // @[cache.scala 68:31]
  wire  _off_T = to_sram_r_ready & to_sram_r_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _off_T_2 = off + 4'h1; // @[cache.scala 69:51]
  wire [3:0] _off_T_3 = _off_T ? _off_T_2 : off; // @[cache.scala 69:31]
  wire [2:0] _GEN_513 = 3'h4 == state_cache ? 3'h1 : state_cache; // @[cache.scala 49:26 74:25 48:30]
  wire [2:0] _GEN_514 = 3'h3 == state_cache ? _state_cache_T_3 : _GEN_513; // @[cache.scala 49:26 68:25]
  wire [3:0] _GEN_515 = 3'h3 == state_cache ? _off_T_3 : off; // @[cache.scala 45:24 49:26 69:25]
  wire  _T_6 = state_cache == 3'h3; // @[cache.scala 80:24]
  wire  _GEN_7184 = 6'h0 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7185 = 4'h0 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7187 = 4'h1 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7189 = 4'h2 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7191 = 4'h3 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7193 = 4'h4 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7195 = 4'h5 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7197 = 4'h6 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7199 = 4'h7 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7201 = 4'h8 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7203 = 4'h9 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7205 = 4'ha == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7207 = 4'hb == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7209 = 4'hc == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7211 = 4'hd == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7213 = 4'he == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7215 = 4'hf == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7216 = 6'h1 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7248 = 6'h2 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7280 = 6'h3 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7312 = 6'h4 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7344 = 6'h5 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7376 = 6'h6 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7408 = 6'h7 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7440 = 6'h8 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7472 = 6'h9 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7504 = 6'ha == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7536 = 6'hb == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7568 = 6'hc == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7600 = 6'hd == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7632 = 6'he == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7664 = 6'hf == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7696 = 6'h10 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7728 = 6'h11 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7760 = 6'h12 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7792 = 6'h13 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7824 = 6'h14 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7856 = 6'h15 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7888 = 6'h16 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7920 = 6'h17 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7952 = 6'h18 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_7984 = 6'h19 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8016 = 6'h1a == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8048 = 6'h1b == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8080 = 6'h1c == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8112 = 6'h1d == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8144 = 6'h1e == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8176 = 6'h1f == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8208 = 6'h20 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8240 = 6'h21 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8272 = 6'h22 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8304 = 6'h23 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8336 = 6'h24 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8368 = 6'h25 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8400 = 6'h26 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8432 = 6'h27 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8464 = 6'h28 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8496 = 6'h29 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8528 = 6'h2a == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8560 = 6'h2b == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8592 = 6'h2c == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8624 = 6'h2d == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8656 = 6'h2e == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8688 = 6'h2f == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8720 = 6'h30 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8752 = 6'h31 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8784 = 6'h32 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8816 = 6'h33 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8848 = 6'h34 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8880 = 6'h35 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8912 = 6'h36 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8944 = 6'h37 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_8976 = 6'h38 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9008 = 6'h39 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9040 = 6'h3a == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9072 = 6'h3b == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9104 = 6'h3c == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9136 = 6'h3d == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9168 = 6'h3e == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9200 = 6'h3f == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_9232 = 2'h0 == replace_set; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2573 = 2'h0 == replace_set & _GEN_7184 | validArray_0_0; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2574 = 2'h0 == replace_set & _GEN_7216 | validArray_0_1; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2575 = 2'h0 == replace_set & _GEN_7248 | validArray_0_2; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2576 = 2'h0 == replace_set & _GEN_7280 | validArray_0_3; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2577 = 2'h0 == replace_set & _GEN_7312 | validArray_0_4; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2578 = 2'h0 == replace_set & _GEN_7344 | validArray_0_5; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2579 = 2'h0 == replace_set & _GEN_7376 | validArray_0_6; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2580 = 2'h0 == replace_set & _GEN_7408 | validArray_0_7; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2581 = 2'h0 == replace_set & _GEN_7440 | validArray_0_8; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2582 = 2'h0 == replace_set & _GEN_7472 | validArray_0_9; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2583 = 2'h0 == replace_set & _GEN_7504 | validArray_0_10; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2584 = 2'h0 == replace_set & _GEN_7536 | validArray_0_11; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2585 = 2'h0 == replace_set & _GEN_7568 | validArray_0_12; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2586 = 2'h0 == replace_set & _GEN_7600 | validArray_0_13; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2587 = 2'h0 == replace_set & _GEN_7632 | validArray_0_14; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2588 = 2'h0 == replace_set & _GEN_7664 | validArray_0_15; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2589 = 2'h0 == replace_set & _GEN_7696 | validArray_0_16; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2590 = 2'h0 == replace_set & _GEN_7728 | validArray_0_17; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2591 = 2'h0 == replace_set & _GEN_7760 | validArray_0_18; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2592 = 2'h0 == replace_set & _GEN_7792 | validArray_0_19; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2593 = 2'h0 == replace_set & _GEN_7824 | validArray_0_20; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2594 = 2'h0 == replace_set & _GEN_7856 | validArray_0_21; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2595 = 2'h0 == replace_set & _GEN_7888 | validArray_0_22; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2596 = 2'h0 == replace_set & _GEN_7920 | validArray_0_23; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2597 = 2'h0 == replace_set & _GEN_7952 | validArray_0_24; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2598 = 2'h0 == replace_set & _GEN_7984 | validArray_0_25; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2599 = 2'h0 == replace_set & _GEN_8016 | validArray_0_26; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2600 = 2'h0 == replace_set & _GEN_8048 | validArray_0_27; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2601 = 2'h0 == replace_set & _GEN_8080 | validArray_0_28; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2602 = 2'h0 == replace_set & _GEN_8112 | validArray_0_29; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2603 = 2'h0 == replace_set & _GEN_8144 | validArray_0_30; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2604 = 2'h0 == replace_set & _GEN_8176 | validArray_0_31; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2605 = 2'h0 == replace_set & _GEN_8208 | validArray_0_32; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2606 = 2'h0 == replace_set & _GEN_8240 | validArray_0_33; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2607 = 2'h0 == replace_set & _GEN_8272 | validArray_0_34; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2608 = 2'h0 == replace_set & _GEN_8304 | validArray_0_35; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2609 = 2'h0 == replace_set & _GEN_8336 | validArray_0_36; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2610 = 2'h0 == replace_set & _GEN_8368 | validArray_0_37; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2611 = 2'h0 == replace_set & _GEN_8400 | validArray_0_38; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2612 = 2'h0 == replace_set & _GEN_8432 | validArray_0_39; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2613 = 2'h0 == replace_set & _GEN_8464 | validArray_0_40; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2614 = 2'h0 == replace_set & _GEN_8496 | validArray_0_41; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2615 = 2'h0 == replace_set & _GEN_8528 | validArray_0_42; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2616 = 2'h0 == replace_set & _GEN_8560 | validArray_0_43; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2617 = 2'h0 == replace_set & _GEN_8592 | validArray_0_44; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2618 = 2'h0 == replace_set & _GEN_8624 | validArray_0_45; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2619 = 2'h0 == replace_set & _GEN_8656 | validArray_0_46; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2620 = 2'h0 == replace_set & _GEN_8688 | validArray_0_47; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2621 = 2'h0 == replace_set & _GEN_8720 | validArray_0_48; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2622 = 2'h0 == replace_set & _GEN_8752 | validArray_0_49; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2623 = 2'h0 == replace_set & _GEN_8784 | validArray_0_50; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2624 = 2'h0 == replace_set & _GEN_8816 | validArray_0_51; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2625 = 2'h0 == replace_set & _GEN_8848 | validArray_0_52; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2626 = 2'h0 == replace_set & _GEN_8880 | validArray_0_53; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2627 = 2'h0 == replace_set & _GEN_8912 | validArray_0_54; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2628 = 2'h0 == replace_set & _GEN_8944 | validArray_0_55; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2629 = 2'h0 == replace_set & _GEN_8976 | validArray_0_56; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2630 = 2'h0 == replace_set & _GEN_9008 | validArray_0_57; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2631 = 2'h0 == replace_set & _GEN_9040 | validArray_0_58; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2632 = 2'h0 == replace_set & _GEN_9072 | validArray_0_59; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2633 = 2'h0 == replace_set & _GEN_9104 | validArray_0_60; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2634 = 2'h0 == replace_set & _GEN_9136 | validArray_0_61; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2635 = 2'h0 == replace_set & _GEN_9168 | validArray_0_62; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2636 = 2'h0 == replace_set & _GEN_9200 | validArray_0_63; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_9424 = 2'h1 == replace_set; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2637 = 2'h1 == replace_set & _GEN_7184 | validArray_1_0; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2638 = 2'h1 == replace_set & _GEN_7216 | validArray_1_1; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2639 = 2'h1 == replace_set & _GEN_7248 | validArray_1_2; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2640 = 2'h1 == replace_set & _GEN_7280 | validArray_1_3; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2641 = 2'h1 == replace_set & _GEN_7312 | validArray_1_4; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2642 = 2'h1 == replace_set & _GEN_7344 | validArray_1_5; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2643 = 2'h1 == replace_set & _GEN_7376 | validArray_1_6; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2644 = 2'h1 == replace_set & _GEN_7408 | validArray_1_7; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2645 = 2'h1 == replace_set & _GEN_7440 | validArray_1_8; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2646 = 2'h1 == replace_set & _GEN_7472 | validArray_1_9; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2647 = 2'h1 == replace_set & _GEN_7504 | validArray_1_10; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2648 = 2'h1 == replace_set & _GEN_7536 | validArray_1_11; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2649 = 2'h1 == replace_set & _GEN_7568 | validArray_1_12; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2650 = 2'h1 == replace_set & _GEN_7600 | validArray_1_13; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2651 = 2'h1 == replace_set & _GEN_7632 | validArray_1_14; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2652 = 2'h1 == replace_set & _GEN_7664 | validArray_1_15; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2653 = 2'h1 == replace_set & _GEN_7696 | validArray_1_16; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2654 = 2'h1 == replace_set & _GEN_7728 | validArray_1_17; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2655 = 2'h1 == replace_set & _GEN_7760 | validArray_1_18; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2656 = 2'h1 == replace_set & _GEN_7792 | validArray_1_19; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2657 = 2'h1 == replace_set & _GEN_7824 | validArray_1_20; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2658 = 2'h1 == replace_set & _GEN_7856 | validArray_1_21; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2659 = 2'h1 == replace_set & _GEN_7888 | validArray_1_22; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2660 = 2'h1 == replace_set & _GEN_7920 | validArray_1_23; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2661 = 2'h1 == replace_set & _GEN_7952 | validArray_1_24; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2662 = 2'h1 == replace_set & _GEN_7984 | validArray_1_25; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2663 = 2'h1 == replace_set & _GEN_8016 | validArray_1_26; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2664 = 2'h1 == replace_set & _GEN_8048 | validArray_1_27; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2665 = 2'h1 == replace_set & _GEN_8080 | validArray_1_28; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2666 = 2'h1 == replace_set & _GEN_8112 | validArray_1_29; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2667 = 2'h1 == replace_set & _GEN_8144 | validArray_1_30; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2668 = 2'h1 == replace_set & _GEN_8176 | validArray_1_31; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2669 = 2'h1 == replace_set & _GEN_8208 | validArray_1_32; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2670 = 2'h1 == replace_set & _GEN_8240 | validArray_1_33; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2671 = 2'h1 == replace_set & _GEN_8272 | validArray_1_34; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2672 = 2'h1 == replace_set & _GEN_8304 | validArray_1_35; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2673 = 2'h1 == replace_set & _GEN_8336 | validArray_1_36; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2674 = 2'h1 == replace_set & _GEN_8368 | validArray_1_37; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2675 = 2'h1 == replace_set & _GEN_8400 | validArray_1_38; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2676 = 2'h1 == replace_set & _GEN_8432 | validArray_1_39; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2677 = 2'h1 == replace_set & _GEN_8464 | validArray_1_40; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2678 = 2'h1 == replace_set & _GEN_8496 | validArray_1_41; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2679 = 2'h1 == replace_set & _GEN_8528 | validArray_1_42; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2680 = 2'h1 == replace_set & _GEN_8560 | validArray_1_43; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2681 = 2'h1 == replace_set & _GEN_8592 | validArray_1_44; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2682 = 2'h1 == replace_set & _GEN_8624 | validArray_1_45; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2683 = 2'h1 == replace_set & _GEN_8656 | validArray_1_46; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2684 = 2'h1 == replace_set & _GEN_8688 | validArray_1_47; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2685 = 2'h1 == replace_set & _GEN_8720 | validArray_1_48; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2686 = 2'h1 == replace_set & _GEN_8752 | validArray_1_49; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2687 = 2'h1 == replace_set & _GEN_8784 | validArray_1_50; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2688 = 2'h1 == replace_set & _GEN_8816 | validArray_1_51; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2689 = 2'h1 == replace_set & _GEN_8848 | validArray_1_52; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2690 = 2'h1 == replace_set & _GEN_8880 | validArray_1_53; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2691 = 2'h1 == replace_set & _GEN_8912 | validArray_1_54; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2692 = 2'h1 == replace_set & _GEN_8944 | validArray_1_55; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2693 = 2'h1 == replace_set & _GEN_8976 | validArray_1_56; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2694 = 2'h1 == replace_set & _GEN_9008 | validArray_1_57; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2695 = 2'h1 == replace_set & _GEN_9040 | validArray_1_58; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2696 = 2'h1 == replace_set & _GEN_9072 | validArray_1_59; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2697 = 2'h1 == replace_set & _GEN_9104 | validArray_1_60; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2698 = 2'h1 == replace_set & _GEN_9136 | validArray_1_61; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2699 = 2'h1 == replace_set & _GEN_9168 | validArray_1_62; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2700 = 2'h1 == replace_set & _GEN_9200 | validArray_1_63; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_9616 = 2'h2 == replace_set; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2701 = 2'h2 == replace_set & _GEN_7184 | validArray_2_0; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2702 = 2'h2 == replace_set & _GEN_7216 | validArray_2_1; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2703 = 2'h2 == replace_set & _GEN_7248 | validArray_2_2; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2704 = 2'h2 == replace_set & _GEN_7280 | validArray_2_3; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2705 = 2'h2 == replace_set & _GEN_7312 | validArray_2_4; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2706 = 2'h2 == replace_set & _GEN_7344 | validArray_2_5; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2707 = 2'h2 == replace_set & _GEN_7376 | validArray_2_6; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2708 = 2'h2 == replace_set & _GEN_7408 | validArray_2_7; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2709 = 2'h2 == replace_set & _GEN_7440 | validArray_2_8; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2710 = 2'h2 == replace_set & _GEN_7472 | validArray_2_9; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2711 = 2'h2 == replace_set & _GEN_7504 | validArray_2_10; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2712 = 2'h2 == replace_set & _GEN_7536 | validArray_2_11; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2713 = 2'h2 == replace_set & _GEN_7568 | validArray_2_12; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2714 = 2'h2 == replace_set & _GEN_7600 | validArray_2_13; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2715 = 2'h2 == replace_set & _GEN_7632 | validArray_2_14; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2716 = 2'h2 == replace_set & _GEN_7664 | validArray_2_15; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2717 = 2'h2 == replace_set & _GEN_7696 | validArray_2_16; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2718 = 2'h2 == replace_set & _GEN_7728 | validArray_2_17; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2719 = 2'h2 == replace_set & _GEN_7760 | validArray_2_18; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2720 = 2'h2 == replace_set & _GEN_7792 | validArray_2_19; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2721 = 2'h2 == replace_set & _GEN_7824 | validArray_2_20; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2722 = 2'h2 == replace_set & _GEN_7856 | validArray_2_21; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2723 = 2'h2 == replace_set & _GEN_7888 | validArray_2_22; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2724 = 2'h2 == replace_set & _GEN_7920 | validArray_2_23; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2725 = 2'h2 == replace_set & _GEN_7952 | validArray_2_24; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2726 = 2'h2 == replace_set & _GEN_7984 | validArray_2_25; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2727 = 2'h2 == replace_set & _GEN_8016 | validArray_2_26; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2728 = 2'h2 == replace_set & _GEN_8048 | validArray_2_27; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2729 = 2'h2 == replace_set & _GEN_8080 | validArray_2_28; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2730 = 2'h2 == replace_set & _GEN_8112 | validArray_2_29; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2731 = 2'h2 == replace_set & _GEN_8144 | validArray_2_30; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2732 = 2'h2 == replace_set & _GEN_8176 | validArray_2_31; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2733 = 2'h2 == replace_set & _GEN_8208 | validArray_2_32; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2734 = 2'h2 == replace_set & _GEN_8240 | validArray_2_33; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2735 = 2'h2 == replace_set & _GEN_8272 | validArray_2_34; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2736 = 2'h2 == replace_set & _GEN_8304 | validArray_2_35; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2737 = 2'h2 == replace_set & _GEN_8336 | validArray_2_36; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2738 = 2'h2 == replace_set & _GEN_8368 | validArray_2_37; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2739 = 2'h2 == replace_set & _GEN_8400 | validArray_2_38; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2740 = 2'h2 == replace_set & _GEN_8432 | validArray_2_39; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2741 = 2'h2 == replace_set & _GEN_8464 | validArray_2_40; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2742 = 2'h2 == replace_set & _GEN_8496 | validArray_2_41; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2743 = 2'h2 == replace_set & _GEN_8528 | validArray_2_42; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2744 = 2'h2 == replace_set & _GEN_8560 | validArray_2_43; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2745 = 2'h2 == replace_set & _GEN_8592 | validArray_2_44; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2746 = 2'h2 == replace_set & _GEN_8624 | validArray_2_45; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2747 = 2'h2 == replace_set & _GEN_8656 | validArray_2_46; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2748 = 2'h2 == replace_set & _GEN_8688 | validArray_2_47; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2749 = 2'h2 == replace_set & _GEN_8720 | validArray_2_48; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2750 = 2'h2 == replace_set & _GEN_8752 | validArray_2_49; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2751 = 2'h2 == replace_set & _GEN_8784 | validArray_2_50; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2752 = 2'h2 == replace_set & _GEN_8816 | validArray_2_51; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2753 = 2'h2 == replace_set & _GEN_8848 | validArray_2_52; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2754 = 2'h2 == replace_set & _GEN_8880 | validArray_2_53; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2755 = 2'h2 == replace_set & _GEN_8912 | validArray_2_54; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2756 = 2'h2 == replace_set & _GEN_8944 | validArray_2_55; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2757 = 2'h2 == replace_set & _GEN_8976 | validArray_2_56; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2758 = 2'h2 == replace_set & _GEN_9008 | validArray_2_57; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2759 = 2'h2 == replace_set & _GEN_9040 | validArray_2_58; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2760 = 2'h2 == replace_set & _GEN_9072 | validArray_2_59; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2761 = 2'h2 == replace_set & _GEN_9104 | validArray_2_60; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2762 = 2'h2 == replace_set & _GEN_9136 | validArray_2_61; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2763 = 2'h2 == replace_set & _GEN_9168 | validArray_2_62; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2764 = 2'h2 == replace_set & _GEN_9200 | validArray_2_63; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_9808 = 2'h3 == replace_set; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2765 = 2'h3 == replace_set & _GEN_7184 | validArray_3_0; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2766 = 2'h3 == replace_set & _GEN_7216 | validArray_3_1; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2767 = 2'h3 == replace_set & _GEN_7248 | validArray_3_2; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2768 = 2'h3 == replace_set & _GEN_7280 | validArray_3_3; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2769 = 2'h3 == replace_set & _GEN_7312 | validArray_3_4; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2770 = 2'h3 == replace_set & _GEN_7344 | validArray_3_5; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2771 = 2'h3 == replace_set & _GEN_7376 | validArray_3_6; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2772 = 2'h3 == replace_set & _GEN_7408 | validArray_3_7; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2773 = 2'h3 == replace_set & _GEN_7440 | validArray_3_8; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2774 = 2'h3 == replace_set & _GEN_7472 | validArray_3_9; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2775 = 2'h3 == replace_set & _GEN_7504 | validArray_3_10; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2776 = 2'h3 == replace_set & _GEN_7536 | validArray_3_11; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2777 = 2'h3 == replace_set & _GEN_7568 | validArray_3_12; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2778 = 2'h3 == replace_set & _GEN_7600 | validArray_3_13; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2779 = 2'h3 == replace_set & _GEN_7632 | validArray_3_14; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2780 = 2'h3 == replace_set & _GEN_7664 | validArray_3_15; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2781 = 2'h3 == replace_set & _GEN_7696 | validArray_3_16; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2782 = 2'h3 == replace_set & _GEN_7728 | validArray_3_17; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2783 = 2'h3 == replace_set & _GEN_7760 | validArray_3_18; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2784 = 2'h3 == replace_set & _GEN_7792 | validArray_3_19; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2785 = 2'h3 == replace_set & _GEN_7824 | validArray_3_20; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2786 = 2'h3 == replace_set & _GEN_7856 | validArray_3_21; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2787 = 2'h3 == replace_set & _GEN_7888 | validArray_3_22; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2788 = 2'h3 == replace_set & _GEN_7920 | validArray_3_23; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2789 = 2'h3 == replace_set & _GEN_7952 | validArray_3_24; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2790 = 2'h3 == replace_set & _GEN_7984 | validArray_3_25; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2791 = 2'h3 == replace_set & _GEN_8016 | validArray_3_26; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2792 = 2'h3 == replace_set & _GEN_8048 | validArray_3_27; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2793 = 2'h3 == replace_set & _GEN_8080 | validArray_3_28; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2794 = 2'h3 == replace_set & _GEN_8112 | validArray_3_29; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2795 = 2'h3 == replace_set & _GEN_8144 | validArray_3_30; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2796 = 2'h3 == replace_set & _GEN_8176 | validArray_3_31; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2797 = 2'h3 == replace_set & _GEN_8208 | validArray_3_32; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2798 = 2'h3 == replace_set & _GEN_8240 | validArray_3_33; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2799 = 2'h3 == replace_set & _GEN_8272 | validArray_3_34; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2800 = 2'h3 == replace_set & _GEN_8304 | validArray_3_35; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2801 = 2'h3 == replace_set & _GEN_8336 | validArray_3_36; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2802 = 2'h3 == replace_set & _GEN_8368 | validArray_3_37; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2803 = 2'h3 == replace_set & _GEN_8400 | validArray_3_38; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2804 = 2'h3 == replace_set & _GEN_8432 | validArray_3_39; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2805 = 2'h3 == replace_set & _GEN_8464 | validArray_3_40; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2806 = 2'h3 == replace_set & _GEN_8496 | validArray_3_41; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2807 = 2'h3 == replace_set & _GEN_8528 | validArray_3_42; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2808 = 2'h3 == replace_set & _GEN_8560 | validArray_3_43; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2809 = 2'h3 == replace_set & _GEN_8592 | validArray_3_44; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2810 = 2'h3 == replace_set & _GEN_8624 | validArray_3_45; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2811 = 2'h3 == replace_set & _GEN_8656 | validArray_3_46; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2812 = 2'h3 == replace_set & _GEN_8688 | validArray_3_47; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2813 = 2'h3 == replace_set & _GEN_8720 | validArray_3_48; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2814 = 2'h3 == replace_set & _GEN_8752 | validArray_3_49; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2815 = 2'h3 == replace_set & _GEN_8784 | validArray_3_50; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2816 = 2'h3 == replace_set & _GEN_8816 | validArray_3_51; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2817 = 2'h3 == replace_set & _GEN_8848 | validArray_3_52; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2818 = 2'h3 == replace_set & _GEN_8880 | validArray_3_53; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2819 = 2'h3 == replace_set & _GEN_8912 | validArray_3_54; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2820 = 2'h3 == replace_set & _GEN_8944 | validArray_3_55; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2821 = 2'h3 == replace_set & _GEN_8976 | validArray_3_56; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2822 = 2'h3 == replace_set & _GEN_9008 | validArray_3_57; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2823 = 2'h3 == replace_set & _GEN_9040 | validArray_3_58; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2824 = 2'h3 == replace_set & _GEN_9072 | validArray_3_59; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2825 = 2'h3 == replace_set & _GEN_9104 | validArray_3_60; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2826 = 2'h3 == replace_set & _GEN_9136 | validArray_3_61; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2827 = 2'h3 == replace_set & _GEN_9168 | validArray_3_62; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_2828 = 2'h3 == replace_set & _GEN_9200 | validArray_3_63; // @[cache.scala 32:29 83:{50,50}]
  wire [31:0] _to_sram_ar_bits_addr_T = {{6'd0}, from_IFU_bits_addr[31:6]}; // @[cache.scala 91:91]
  wire [37:0] _GEN_10513 = {_to_sram_ar_bits_addr_T, 6'h0}; // @[cache.scala 91:104]
  wire [38:0] _to_sram_ar_bits_addr_T_1 = {{1'd0}, _GEN_10513}; // @[cache.scala 91:104]
  wire [38:0] _to_sram_ar_bits_addr_T_3 = _T_3 ? _to_sram_ar_bits_addr_T_1 : 39'h0; // @[Mux.scala 81:58]
  wire [3:0] _to_sram_ar_bits_len_T_1 = _T_3 ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [31:0] _GEN_6160 = dataArray_0_0_cachedata_MPORT_data; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6161 = _GEN_7184 & 4'h1 == EntId[3:0] ? dataArray_0_1_cachedata_MPORT_data : _GEN_6160; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6162 = _GEN_7184 & 4'h2 == EntId[3:0] ? dataArray_0_2_cachedata_MPORT_data : _GEN_6161; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6163 = _GEN_7184 & 4'h3 == EntId[3:0] ? dataArray_0_3_cachedata_MPORT_data : _GEN_6162; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6164 = _GEN_7184 & 4'h4 == EntId[3:0] ? dataArray_0_4_cachedata_MPORT_data : _GEN_6163; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6165 = _GEN_7184 & 4'h5 == EntId[3:0] ? dataArray_0_5_cachedata_MPORT_data : _GEN_6164; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6166 = _GEN_7184 & 4'h6 == EntId[3:0] ? dataArray_0_6_cachedata_MPORT_data : _GEN_6165; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6167 = _GEN_7184 & 4'h7 == EntId[3:0] ? dataArray_0_7_cachedata_MPORT_data : _GEN_6166; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6168 = _GEN_7184 & 4'h8 == EntId[3:0] ? dataArray_0_8_cachedata_MPORT_data : _GEN_6167; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6169 = _GEN_7184 & 4'h9 == EntId[3:0] ? dataArray_0_9_cachedata_MPORT_data : _GEN_6168; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6170 = _GEN_7184 & 4'ha == EntId[3:0] ? dataArray_0_10_cachedata_MPORT_data : _GEN_6169; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6171 = _GEN_7184 & 4'hb == EntId[3:0] ? dataArray_0_11_cachedata_MPORT_data : _GEN_6170; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6172 = _GEN_7184 & 4'hc == EntId[3:0] ? dataArray_0_12_cachedata_MPORT_data : _GEN_6171; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6173 = _GEN_7184 & 4'hd == EntId[3:0] ? dataArray_0_13_cachedata_MPORT_data : _GEN_6172; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6174 = _GEN_7184 & 4'he == EntId[3:0] ? dataArray_0_14_cachedata_MPORT_data : _GEN_6173; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6175 = _GEN_7184 & 4'hf == EntId[3:0] ? dataArray_0_15_cachedata_MPORT_data : _GEN_6174; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6176 = _GEN_7216 & 4'h0 == EntId[3:0] ? dataArray_1_0_cachedata_MPORT_data : _GEN_6175; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6177 = _GEN_7216 & 4'h1 == EntId[3:0] ? dataArray_1_1_cachedata_MPORT_data : _GEN_6176; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6178 = _GEN_7216 & 4'h2 == EntId[3:0] ? dataArray_1_2_cachedata_MPORT_data : _GEN_6177; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6179 = _GEN_7216 & 4'h3 == EntId[3:0] ? dataArray_1_3_cachedata_MPORT_data : _GEN_6178; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6180 = _GEN_7216 & 4'h4 == EntId[3:0] ? dataArray_1_4_cachedata_MPORT_data : _GEN_6179; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6181 = _GEN_7216 & 4'h5 == EntId[3:0] ? dataArray_1_5_cachedata_MPORT_data : _GEN_6180; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6182 = _GEN_7216 & 4'h6 == EntId[3:0] ? dataArray_1_6_cachedata_MPORT_data : _GEN_6181; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6183 = _GEN_7216 & 4'h7 == EntId[3:0] ? dataArray_1_7_cachedata_MPORT_data : _GEN_6182; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6184 = _GEN_7216 & 4'h8 == EntId[3:0] ? dataArray_1_8_cachedata_MPORT_data : _GEN_6183; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6185 = _GEN_7216 & 4'h9 == EntId[3:0] ? dataArray_1_9_cachedata_MPORT_data : _GEN_6184; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6186 = _GEN_7216 & 4'ha == EntId[3:0] ? dataArray_1_10_cachedata_MPORT_data : _GEN_6185; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6187 = _GEN_7216 & 4'hb == EntId[3:0] ? dataArray_1_11_cachedata_MPORT_data : _GEN_6186; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6188 = _GEN_7216 & 4'hc == EntId[3:0] ? dataArray_1_12_cachedata_MPORT_data : _GEN_6187; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6189 = _GEN_7216 & 4'hd == EntId[3:0] ? dataArray_1_13_cachedata_MPORT_data : _GEN_6188; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6190 = _GEN_7216 & 4'he == EntId[3:0] ? dataArray_1_14_cachedata_MPORT_data : _GEN_6189; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6191 = _GEN_7216 & 4'hf == EntId[3:0] ? dataArray_1_15_cachedata_MPORT_data : _GEN_6190; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6192 = _GEN_7248 & 4'h0 == EntId[3:0] ? dataArray_2_0_cachedata_MPORT_data : _GEN_6191; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6193 = _GEN_7248 & 4'h1 == EntId[3:0] ? dataArray_2_1_cachedata_MPORT_data : _GEN_6192; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6194 = _GEN_7248 & 4'h2 == EntId[3:0] ? dataArray_2_2_cachedata_MPORT_data : _GEN_6193; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6195 = _GEN_7248 & 4'h3 == EntId[3:0] ? dataArray_2_3_cachedata_MPORT_data : _GEN_6194; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6196 = _GEN_7248 & 4'h4 == EntId[3:0] ? dataArray_2_4_cachedata_MPORT_data : _GEN_6195; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6197 = _GEN_7248 & 4'h5 == EntId[3:0] ? dataArray_2_5_cachedata_MPORT_data : _GEN_6196; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6198 = _GEN_7248 & 4'h6 == EntId[3:0] ? dataArray_2_6_cachedata_MPORT_data : _GEN_6197; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6199 = _GEN_7248 & 4'h7 == EntId[3:0] ? dataArray_2_7_cachedata_MPORT_data : _GEN_6198; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6200 = _GEN_7248 & 4'h8 == EntId[3:0] ? dataArray_2_8_cachedata_MPORT_data : _GEN_6199; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6201 = _GEN_7248 & 4'h9 == EntId[3:0] ? dataArray_2_9_cachedata_MPORT_data : _GEN_6200; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6202 = _GEN_7248 & 4'ha == EntId[3:0] ? dataArray_2_10_cachedata_MPORT_data : _GEN_6201; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6203 = _GEN_7248 & 4'hb == EntId[3:0] ? dataArray_2_11_cachedata_MPORT_data : _GEN_6202; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6204 = _GEN_7248 & 4'hc == EntId[3:0] ? dataArray_2_12_cachedata_MPORT_data : _GEN_6203; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6205 = _GEN_7248 & 4'hd == EntId[3:0] ? dataArray_2_13_cachedata_MPORT_data : _GEN_6204; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6206 = _GEN_7248 & 4'he == EntId[3:0] ? dataArray_2_14_cachedata_MPORT_data : _GEN_6205; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6207 = _GEN_7248 & 4'hf == EntId[3:0] ? dataArray_2_15_cachedata_MPORT_data : _GEN_6206; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6208 = _GEN_7280 & 4'h0 == EntId[3:0] ? dataArray_3_0_cachedata_MPORT_data : _GEN_6207; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6209 = _GEN_7280 & 4'h1 == EntId[3:0] ? dataArray_3_1_cachedata_MPORT_data : _GEN_6208; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6210 = _GEN_7280 & 4'h2 == EntId[3:0] ? dataArray_3_2_cachedata_MPORT_data : _GEN_6209; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6211 = _GEN_7280 & 4'h3 == EntId[3:0] ? dataArray_3_3_cachedata_MPORT_data : _GEN_6210; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6212 = _GEN_7280 & 4'h4 == EntId[3:0] ? dataArray_3_4_cachedata_MPORT_data : _GEN_6211; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6213 = _GEN_7280 & 4'h5 == EntId[3:0] ? dataArray_3_5_cachedata_MPORT_data : _GEN_6212; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6214 = _GEN_7280 & 4'h6 == EntId[3:0] ? dataArray_3_6_cachedata_MPORT_data : _GEN_6213; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6215 = _GEN_7280 & 4'h7 == EntId[3:0] ? dataArray_3_7_cachedata_MPORT_data : _GEN_6214; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6216 = _GEN_7280 & 4'h8 == EntId[3:0] ? dataArray_3_8_cachedata_MPORT_data : _GEN_6215; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6217 = _GEN_7280 & 4'h9 == EntId[3:0] ? dataArray_3_9_cachedata_MPORT_data : _GEN_6216; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6218 = _GEN_7280 & 4'ha == EntId[3:0] ? dataArray_3_10_cachedata_MPORT_data : _GEN_6217; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6219 = _GEN_7280 & 4'hb == EntId[3:0] ? dataArray_3_11_cachedata_MPORT_data : _GEN_6218; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6220 = _GEN_7280 & 4'hc == EntId[3:0] ? dataArray_3_12_cachedata_MPORT_data : _GEN_6219; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6221 = _GEN_7280 & 4'hd == EntId[3:0] ? dataArray_3_13_cachedata_MPORT_data : _GEN_6220; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6222 = _GEN_7280 & 4'he == EntId[3:0] ? dataArray_3_14_cachedata_MPORT_data : _GEN_6221; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6223 = _GEN_7280 & 4'hf == EntId[3:0] ? dataArray_3_15_cachedata_MPORT_data : _GEN_6222; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6224 = _GEN_7312 & 4'h0 == EntId[3:0] ? dataArray_4_0_cachedata_MPORT_data : _GEN_6223; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6225 = _GEN_7312 & 4'h1 == EntId[3:0] ? dataArray_4_1_cachedata_MPORT_data : _GEN_6224; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6226 = _GEN_7312 & 4'h2 == EntId[3:0] ? dataArray_4_2_cachedata_MPORT_data : _GEN_6225; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6227 = _GEN_7312 & 4'h3 == EntId[3:0] ? dataArray_4_3_cachedata_MPORT_data : _GEN_6226; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6228 = _GEN_7312 & 4'h4 == EntId[3:0] ? dataArray_4_4_cachedata_MPORT_data : _GEN_6227; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6229 = _GEN_7312 & 4'h5 == EntId[3:0] ? dataArray_4_5_cachedata_MPORT_data : _GEN_6228; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6230 = _GEN_7312 & 4'h6 == EntId[3:0] ? dataArray_4_6_cachedata_MPORT_data : _GEN_6229; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6231 = _GEN_7312 & 4'h7 == EntId[3:0] ? dataArray_4_7_cachedata_MPORT_data : _GEN_6230; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6232 = _GEN_7312 & 4'h8 == EntId[3:0] ? dataArray_4_8_cachedata_MPORT_data : _GEN_6231; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6233 = _GEN_7312 & 4'h9 == EntId[3:0] ? dataArray_4_9_cachedata_MPORT_data : _GEN_6232; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6234 = _GEN_7312 & 4'ha == EntId[3:0] ? dataArray_4_10_cachedata_MPORT_data : _GEN_6233; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6235 = _GEN_7312 & 4'hb == EntId[3:0] ? dataArray_4_11_cachedata_MPORT_data : _GEN_6234; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6236 = _GEN_7312 & 4'hc == EntId[3:0] ? dataArray_4_12_cachedata_MPORT_data : _GEN_6235; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6237 = _GEN_7312 & 4'hd == EntId[3:0] ? dataArray_4_13_cachedata_MPORT_data : _GEN_6236; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6238 = _GEN_7312 & 4'he == EntId[3:0] ? dataArray_4_14_cachedata_MPORT_data : _GEN_6237; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6239 = _GEN_7312 & 4'hf == EntId[3:0] ? dataArray_4_15_cachedata_MPORT_data : _GEN_6238; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6240 = _GEN_7344 & 4'h0 == EntId[3:0] ? dataArray_5_0_cachedata_MPORT_data : _GEN_6239; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6241 = _GEN_7344 & 4'h1 == EntId[3:0] ? dataArray_5_1_cachedata_MPORT_data : _GEN_6240; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6242 = _GEN_7344 & 4'h2 == EntId[3:0] ? dataArray_5_2_cachedata_MPORT_data : _GEN_6241; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6243 = _GEN_7344 & 4'h3 == EntId[3:0] ? dataArray_5_3_cachedata_MPORT_data : _GEN_6242; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6244 = _GEN_7344 & 4'h4 == EntId[3:0] ? dataArray_5_4_cachedata_MPORT_data : _GEN_6243; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6245 = _GEN_7344 & 4'h5 == EntId[3:0] ? dataArray_5_5_cachedata_MPORT_data : _GEN_6244; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6246 = _GEN_7344 & 4'h6 == EntId[3:0] ? dataArray_5_6_cachedata_MPORT_data : _GEN_6245; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6247 = _GEN_7344 & 4'h7 == EntId[3:0] ? dataArray_5_7_cachedata_MPORT_data : _GEN_6246; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6248 = _GEN_7344 & 4'h8 == EntId[3:0] ? dataArray_5_8_cachedata_MPORT_data : _GEN_6247; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6249 = _GEN_7344 & 4'h9 == EntId[3:0] ? dataArray_5_9_cachedata_MPORT_data : _GEN_6248; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6250 = _GEN_7344 & 4'ha == EntId[3:0] ? dataArray_5_10_cachedata_MPORT_data : _GEN_6249; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6251 = _GEN_7344 & 4'hb == EntId[3:0] ? dataArray_5_11_cachedata_MPORT_data : _GEN_6250; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6252 = _GEN_7344 & 4'hc == EntId[3:0] ? dataArray_5_12_cachedata_MPORT_data : _GEN_6251; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6253 = _GEN_7344 & 4'hd == EntId[3:0] ? dataArray_5_13_cachedata_MPORT_data : _GEN_6252; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6254 = _GEN_7344 & 4'he == EntId[3:0] ? dataArray_5_14_cachedata_MPORT_data : _GEN_6253; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6255 = _GEN_7344 & 4'hf == EntId[3:0] ? dataArray_5_15_cachedata_MPORT_data : _GEN_6254; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6256 = _GEN_7376 & 4'h0 == EntId[3:0] ? dataArray_6_0_cachedata_MPORT_data : _GEN_6255; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6257 = _GEN_7376 & 4'h1 == EntId[3:0] ? dataArray_6_1_cachedata_MPORT_data : _GEN_6256; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6258 = _GEN_7376 & 4'h2 == EntId[3:0] ? dataArray_6_2_cachedata_MPORT_data : _GEN_6257; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6259 = _GEN_7376 & 4'h3 == EntId[3:0] ? dataArray_6_3_cachedata_MPORT_data : _GEN_6258; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6260 = _GEN_7376 & 4'h4 == EntId[3:0] ? dataArray_6_4_cachedata_MPORT_data : _GEN_6259; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6261 = _GEN_7376 & 4'h5 == EntId[3:0] ? dataArray_6_5_cachedata_MPORT_data : _GEN_6260; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6262 = _GEN_7376 & 4'h6 == EntId[3:0] ? dataArray_6_6_cachedata_MPORT_data : _GEN_6261; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6263 = _GEN_7376 & 4'h7 == EntId[3:0] ? dataArray_6_7_cachedata_MPORT_data : _GEN_6262; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6264 = _GEN_7376 & 4'h8 == EntId[3:0] ? dataArray_6_8_cachedata_MPORT_data : _GEN_6263; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6265 = _GEN_7376 & 4'h9 == EntId[3:0] ? dataArray_6_9_cachedata_MPORT_data : _GEN_6264; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6266 = _GEN_7376 & 4'ha == EntId[3:0] ? dataArray_6_10_cachedata_MPORT_data : _GEN_6265; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6267 = _GEN_7376 & 4'hb == EntId[3:0] ? dataArray_6_11_cachedata_MPORT_data : _GEN_6266; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6268 = _GEN_7376 & 4'hc == EntId[3:0] ? dataArray_6_12_cachedata_MPORT_data : _GEN_6267; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6269 = _GEN_7376 & 4'hd == EntId[3:0] ? dataArray_6_13_cachedata_MPORT_data : _GEN_6268; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6270 = _GEN_7376 & 4'he == EntId[3:0] ? dataArray_6_14_cachedata_MPORT_data : _GEN_6269; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6271 = _GEN_7376 & 4'hf == EntId[3:0] ? dataArray_6_15_cachedata_MPORT_data : _GEN_6270; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6272 = _GEN_7408 & 4'h0 == EntId[3:0] ? dataArray_7_0_cachedata_MPORT_data : _GEN_6271; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6273 = _GEN_7408 & 4'h1 == EntId[3:0] ? dataArray_7_1_cachedata_MPORT_data : _GEN_6272; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6274 = _GEN_7408 & 4'h2 == EntId[3:0] ? dataArray_7_2_cachedata_MPORT_data : _GEN_6273; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6275 = _GEN_7408 & 4'h3 == EntId[3:0] ? dataArray_7_3_cachedata_MPORT_data : _GEN_6274; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6276 = _GEN_7408 & 4'h4 == EntId[3:0] ? dataArray_7_4_cachedata_MPORT_data : _GEN_6275; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6277 = _GEN_7408 & 4'h5 == EntId[3:0] ? dataArray_7_5_cachedata_MPORT_data : _GEN_6276; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6278 = _GEN_7408 & 4'h6 == EntId[3:0] ? dataArray_7_6_cachedata_MPORT_data : _GEN_6277; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6279 = _GEN_7408 & 4'h7 == EntId[3:0] ? dataArray_7_7_cachedata_MPORT_data : _GEN_6278; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6280 = _GEN_7408 & 4'h8 == EntId[3:0] ? dataArray_7_8_cachedata_MPORT_data : _GEN_6279; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6281 = _GEN_7408 & 4'h9 == EntId[3:0] ? dataArray_7_9_cachedata_MPORT_data : _GEN_6280; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6282 = _GEN_7408 & 4'ha == EntId[3:0] ? dataArray_7_10_cachedata_MPORT_data : _GEN_6281; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6283 = _GEN_7408 & 4'hb == EntId[3:0] ? dataArray_7_11_cachedata_MPORT_data : _GEN_6282; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6284 = _GEN_7408 & 4'hc == EntId[3:0] ? dataArray_7_12_cachedata_MPORT_data : _GEN_6283; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6285 = _GEN_7408 & 4'hd == EntId[3:0] ? dataArray_7_13_cachedata_MPORT_data : _GEN_6284; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6286 = _GEN_7408 & 4'he == EntId[3:0] ? dataArray_7_14_cachedata_MPORT_data : _GEN_6285; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6287 = _GEN_7408 & 4'hf == EntId[3:0] ? dataArray_7_15_cachedata_MPORT_data : _GEN_6286; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6288 = _GEN_7440 & 4'h0 == EntId[3:0] ? dataArray_8_0_cachedata_MPORT_data : _GEN_6287; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6289 = _GEN_7440 & 4'h1 == EntId[3:0] ? dataArray_8_1_cachedata_MPORT_data : _GEN_6288; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6290 = _GEN_7440 & 4'h2 == EntId[3:0] ? dataArray_8_2_cachedata_MPORT_data : _GEN_6289; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6291 = _GEN_7440 & 4'h3 == EntId[3:0] ? dataArray_8_3_cachedata_MPORT_data : _GEN_6290; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6292 = _GEN_7440 & 4'h4 == EntId[3:0] ? dataArray_8_4_cachedata_MPORT_data : _GEN_6291; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6293 = _GEN_7440 & 4'h5 == EntId[3:0] ? dataArray_8_5_cachedata_MPORT_data : _GEN_6292; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6294 = _GEN_7440 & 4'h6 == EntId[3:0] ? dataArray_8_6_cachedata_MPORT_data : _GEN_6293; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6295 = _GEN_7440 & 4'h7 == EntId[3:0] ? dataArray_8_7_cachedata_MPORT_data : _GEN_6294; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6296 = _GEN_7440 & 4'h8 == EntId[3:0] ? dataArray_8_8_cachedata_MPORT_data : _GEN_6295; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6297 = _GEN_7440 & 4'h9 == EntId[3:0] ? dataArray_8_9_cachedata_MPORT_data : _GEN_6296; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6298 = _GEN_7440 & 4'ha == EntId[3:0] ? dataArray_8_10_cachedata_MPORT_data : _GEN_6297; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6299 = _GEN_7440 & 4'hb == EntId[3:0] ? dataArray_8_11_cachedata_MPORT_data : _GEN_6298; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6300 = _GEN_7440 & 4'hc == EntId[3:0] ? dataArray_8_12_cachedata_MPORT_data : _GEN_6299; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6301 = _GEN_7440 & 4'hd == EntId[3:0] ? dataArray_8_13_cachedata_MPORT_data : _GEN_6300; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6302 = _GEN_7440 & 4'he == EntId[3:0] ? dataArray_8_14_cachedata_MPORT_data : _GEN_6301; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6303 = _GEN_7440 & 4'hf == EntId[3:0] ? dataArray_8_15_cachedata_MPORT_data : _GEN_6302; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6304 = _GEN_7472 & 4'h0 == EntId[3:0] ? dataArray_9_0_cachedata_MPORT_data : _GEN_6303; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6305 = _GEN_7472 & 4'h1 == EntId[3:0] ? dataArray_9_1_cachedata_MPORT_data : _GEN_6304; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6306 = _GEN_7472 & 4'h2 == EntId[3:0] ? dataArray_9_2_cachedata_MPORT_data : _GEN_6305; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6307 = _GEN_7472 & 4'h3 == EntId[3:0] ? dataArray_9_3_cachedata_MPORT_data : _GEN_6306; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6308 = _GEN_7472 & 4'h4 == EntId[3:0] ? dataArray_9_4_cachedata_MPORT_data : _GEN_6307; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6309 = _GEN_7472 & 4'h5 == EntId[3:0] ? dataArray_9_5_cachedata_MPORT_data : _GEN_6308; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6310 = _GEN_7472 & 4'h6 == EntId[3:0] ? dataArray_9_6_cachedata_MPORT_data : _GEN_6309; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6311 = _GEN_7472 & 4'h7 == EntId[3:0] ? dataArray_9_7_cachedata_MPORT_data : _GEN_6310; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6312 = _GEN_7472 & 4'h8 == EntId[3:0] ? dataArray_9_8_cachedata_MPORT_data : _GEN_6311; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6313 = _GEN_7472 & 4'h9 == EntId[3:0] ? dataArray_9_9_cachedata_MPORT_data : _GEN_6312; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6314 = _GEN_7472 & 4'ha == EntId[3:0] ? dataArray_9_10_cachedata_MPORT_data : _GEN_6313; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6315 = _GEN_7472 & 4'hb == EntId[3:0] ? dataArray_9_11_cachedata_MPORT_data : _GEN_6314; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6316 = _GEN_7472 & 4'hc == EntId[3:0] ? dataArray_9_12_cachedata_MPORT_data : _GEN_6315; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6317 = _GEN_7472 & 4'hd == EntId[3:0] ? dataArray_9_13_cachedata_MPORT_data : _GEN_6316; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6318 = _GEN_7472 & 4'he == EntId[3:0] ? dataArray_9_14_cachedata_MPORT_data : _GEN_6317; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6319 = _GEN_7472 & 4'hf == EntId[3:0] ? dataArray_9_15_cachedata_MPORT_data : _GEN_6318; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6320 = _GEN_7504 & 4'h0 == EntId[3:0] ? dataArray_10_0_cachedata_MPORT_data : _GEN_6319; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6321 = _GEN_7504 & 4'h1 == EntId[3:0] ? dataArray_10_1_cachedata_MPORT_data : _GEN_6320; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6322 = _GEN_7504 & 4'h2 == EntId[3:0] ? dataArray_10_2_cachedata_MPORT_data : _GEN_6321; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6323 = _GEN_7504 & 4'h3 == EntId[3:0] ? dataArray_10_3_cachedata_MPORT_data : _GEN_6322; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6324 = _GEN_7504 & 4'h4 == EntId[3:0] ? dataArray_10_4_cachedata_MPORT_data : _GEN_6323; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6325 = _GEN_7504 & 4'h5 == EntId[3:0] ? dataArray_10_5_cachedata_MPORT_data : _GEN_6324; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6326 = _GEN_7504 & 4'h6 == EntId[3:0] ? dataArray_10_6_cachedata_MPORT_data : _GEN_6325; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6327 = _GEN_7504 & 4'h7 == EntId[3:0] ? dataArray_10_7_cachedata_MPORT_data : _GEN_6326; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6328 = _GEN_7504 & 4'h8 == EntId[3:0] ? dataArray_10_8_cachedata_MPORT_data : _GEN_6327; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6329 = _GEN_7504 & 4'h9 == EntId[3:0] ? dataArray_10_9_cachedata_MPORT_data : _GEN_6328; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6330 = _GEN_7504 & 4'ha == EntId[3:0] ? dataArray_10_10_cachedata_MPORT_data : _GEN_6329; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6331 = _GEN_7504 & 4'hb == EntId[3:0] ? dataArray_10_11_cachedata_MPORT_data : _GEN_6330; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6332 = _GEN_7504 & 4'hc == EntId[3:0] ? dataArray_10_12_cachedata_MPORT_data : _GEN_6331; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6333 = _GEN_7504 & 4'hd == EntId[3:0] ? dataArray_10_13_cachedata_MPORT_data : _GEN_6332; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6334 = _GEN_7504 & 4'he == EntId[3:0] ? dataArray_10_14_cachedata_MPORT_data : _GEN_6333; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6335 = _GEN_7504 & 4'hf == EntId[3:0] ? dataArray_10_15_cachedata_MPORT_data : _GEN_6334; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6336 = _GEN_7536 & 4'h0 == EntId[3:0] ? dataArray_11_0_cachedata_MPORT_data : _GEN_6335; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6337 = _GEN_7536 & 4'h1 == EntId[3:0] ? dataArray_11_1_cachedata_MPORT_data : _GEN_6336; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6338 = _GEN_7536 & 4'h2 == EntId[3:0] ? dataArray_11_2_cachedata_MPORT_data : _GEN_6337; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6339 = _GEN_7536 & 4'h3 == EntId[3:0] ? dataArray_11_3_cachedata_MPORT_data : _GEN_6338; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6340 = _GEN_7536 & 4'h4 == EntId[3:0] ? dataArray_11_4_cachedata_MPORT_data : _GEN_6339; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6341 = _GEN_7536 & 4'h5 == EntId[3:0] ? dataArray_11_5_cachedata_MPORT_data : _GEN_6340; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6342 = _GEN_7536 & 4'h6 == EntId[3:0] ? dataArray_11_6_cachedata_MPORT_data : _GEN_6341; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6343 = _GEN_7536 & 4'h7 == EntId[3:0] ? dataArray_11_7_cachedata_MPORT_data : _GEN_6342; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6344 = _GEN_7536 & 4'h8 == EntId[3:0] ? dataArray_11_8_cachedata_MPORT_data : _GEN_6343; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6345 = _GEN_7536 & 4'h9 == EntId[3:0] ? dataArray_11_9_cachedata_MPORT_data : _GEN_6344; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6346 = _GEN_7536 & 4'ha == EntId[3:0] ? dataArray_11_10_cachedata_MPORT_data : _GEN_6345; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6347 = _GEN_7536 & 4'hb == EntId[3:0] ? dataArray_11_11_cachedata_MPORT_data : _GEN_6346; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6348 = _GEN_7536 & 4'hc == EntId[3:0] ? dataArray_11_12_cachedata_MPORT_data : _GEN_6347; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6349 = _GEN_7536 & 4'hd == EntId[3:0] ? dataArray_11_13_cachedata_MPORT_data : _GEN_6348; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6350 = _GEN_7536 & 4'he == EntId[3:0] ? dataArray_11_14_cachedata_MPORT_data : _GEN_6349; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6351 = _GEN_7536 & 4'hf == EntId[3:0] ? dataArray_11_15_cachedata_MPORT_data : _GEN_6350; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6352 = _GEN_7568 & 4'h0 == EntId[3:0] ? dataArray_12_0_cachedata_MPORT_data : _GEN_6351; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6353 = _GEN_7568 & 4'h1 == EntId[3:0] ? dataArray_12_1_cachedata_MPORT_data : _GEN_6352; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6354 = _GEN_7568 & 4'h2 == EntId[3:0] ? dataArray_12_2_cachedata_MPORT_data : _GEN_6353; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6355 = _GEN_7568 & 4'h3 == EntId[3:0] ? dataArray_12_3_cachedata_MPORT_data : _GEN_6354; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6356 = _GEN_7568 & 4'h4 == EntId[3:0] ? dataArray_12_4_cachedata_MPORT_data : _GEN_6355; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6357 = _GEN_7568 & 4'h5 == EntId[3:0] ? dataArray_12_5_cachedata_MPORT_data : _GEN_6356; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6358 = _GEN_7568 & 4'h6 == EntId[3:0] ? dataArray_12_6_cachedata_MPORT_data : _GEN_6357; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6359 = _GEN_7568 & 4'h7 == EntId[3:0] ? dataArray_12_7_cachedata_MPORT_data : _GEN_6358; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6360 = _GEN_7568 & 4'h8 == EntId[3:0] ? dataArray_12_8_cachedata_MPORT_data : _GEN_6359; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6361 = _GEN_7568 & 4'h9 == EntId[3:0] ? dataArray_12_9_cachedata_MPORT_data : _GEN_6360; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6362 = _GEN_7568 & 4'ha == EntId[3:0] ? dataArray_12_10_cachedata_MPORT_data : _GEN_6361; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6363 = _GEN_7568 & 4'hb == EntId[3:0] ? dataArray_12_11_cachedata_MPORT_data : _GEN_6362; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6364 = _GEN_7568 & 4'hc == EntId[3:0] ? dataArray_12_12_cachedata_MPORT_data : _GEN_6363; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6365 = _GEN_7568 & 4'hd == EntId[3:0] ? dataArray_12_13_cachedata_MPORT_data : _GEN_6364; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6366 = _GEN_7568 & 4'he == EntId[3:0] ? dataArray_12_14_cachedata_MPORT_data : _GEN_6365; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6367 = _GEN_7568 & 4'hf == EntId[3:0] ? dataArray_12_15_cachedata_MPORT_data : _GEN_6366; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6368 = _GEN_7600 & 4'h0 == EntId[3:0] ? dataArray_13_0_cachedata_MPORT_data : _GEN_6367; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6369 = _GEN_7600 & 4'h1 == EntId[3:0] ? dataArray_13_1_cachedata_MPORT_data : _GEN_6368; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6370 = _GEN_7600 & 4'h2 == EntId[3:0] ? dataArray_13_2_cachedata_MPORT_data : _GEN_6369; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6371 = _GEN_7600 & 4'h3 == EntId[3:0] ? dataArray_13_3_cachedata_MPORT_data : _GEN_6370; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6372 = _GEN_7600 & 4'h4 == EntId[3:0] ? dataArray_13_4_cachedata_MPORT_data : _GEN_6371; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6373 = _GEN_7600 & 4'h5 == EntId[3:0] ? dataArray_13_5_cachedata_MPORT_data : _GEN_6372; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6374 = _GEN_7600 & 4'h6 == EntId[3:0] ? dataArray_13_6_cachedata_MPORT_data : _GEN_6373; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6375 = _GEN_7600 & 4'h7 == EntId[3:0] ? dataArray_13_7_cachedata_MPORT_data : _GEN_6374; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6376 = _GEN_7600 & 4'h8 == EntId[3:0] ? dataArray_13_8_cachedata_MPORT_data : _GEN_6375; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6377 = _GEN_7600 & 4'h9 == EntId[3:0] ? dataArray_13_9_cachedata_MPORT_data : _GEN_6376; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6378 = _GEN_7600 & 4'ha == EntId[3:0] ? dataArray_13_10_cachedata_MPORT_data : _GEN_6377; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6379 = _GEN_7600 & 4'hb == EntId[3:0] ? dataArray_13_11_cachedata_MPORT_data : _GEN_6378; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6380 = _GEN_7600 & 4'hc == EntId[3:0] ? dataArray_13_12_cachedata_MPORT_data : _GEN_6379; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6381 = _GEN_7600 & 4'hd == EntId[3:0] ? dataArray_13_13_cachedata_MPORT_data : _GEN_6380; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6382 = _GEN_7600 & 4'he == EntId[3:0] ? dataArray_13_14_cachedata_MPORT_data : _GEN_6381; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6383 = _GEN_7600 & 4'hf == EntId[3:0] ? dataArray_13_15_cachedata_MPORT_data : _GEN_6382; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6384 = _GEN_7632 & 4'h0 == EntId[3:0] ? dataArray_14_0_cachedata_MPORT_data : _GEN_6383; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6385 = _GEN_7632 & 4'h1 == EntId[3:0] ? dataArray_14_1_cachedata_MPORT_data : _GEN_6384; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6386 = _GEN_7632 & 4'h2 == EntId[3:0] ? dataArray_14_2_cachedata_MPORT_data : _GEN_6385; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6387 = _GEN_7632 & 4'h3 == EntId[3:0] ? dataArray_14_3_cachedata_MPORT_data : _GEN_6386; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6388 = _GEN_7632 & 4'h4 == EntId[3:0] ? dataArray_14_4_cachedata_MPORT_data : _GEN_6387; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6389 = _GEN_7632 & 4'h5 == EntId[3:0] ? dataArray_14_5_cachedata_MPORT_data : _GEN_6388; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6390 = _GEN_7632 & 4'h6 == EntId[3:0] ? dataArray_14_6_cachedata_MPORT_data : _GEN_6389; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6391 = _GEN_7632 & 4'h7 == EntId[3:0] ? dataArray_14_7_cachedata_MPORT_data : _GEN_6390; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6392 = _GEN_7632 & 4'h8 == EntId[3:0] ? dataArray_14_8_cachedata_MPORT_data : _GEN_6391; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6393 = _GEN_7632 & 4'h9 == EntId[3:0] ? dataArray_14_9_cachedata_MPORT_data : _GEN_6392; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6394 = _GEN_7632 & 4'ha == EntId[3:0] ? dataArray_14_10_cachedata_MPORT_data : _GEN_6393; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6395 = _GEN_7632 & 4'hb == EntId[3:0] ? dataArray_14_11_cachedata_MPORT_data : _GEN_6394; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6396 = _GEN_7632 & 4'hc == EntId[3:0] ? dataArray_14_12_cachedata_MPORT_data : _GEN_6395; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6397 = _GEN_7632 & 4'hd == EntId[3:0] ? dataArray_14_13_cachedata_MPORT_data : _GEN_6396; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6398 = _GEN_7632 & 4'he == EntId[3:0] ? dataArray_14_14_cachedata_MPORT_data : _GEN_6397; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6399 = _GEN_7632 & 4'hf == EntId[3:0] ? dataArray_14_15_cachedata_MPORT_data : _GEN_6398; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6400 = _GEN_7664 & 4'h0 == EntId[3:0] ? dataArray_15_0_cachedata_MPORT_data : _GEN_6399; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6401 = _GEN_7664 & 4'h1 == EntId[3:0] ? dataArray_15_1_cachedata_MPORT_data : _GEN_6400; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6402 = _GEN_7664 & 4'h2 == EntId[3:0] ? dataArray_15_2_cachedata_MPORT_data : _GEN_6401; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6403 = _GEN_7664 & 4'h3 == EntId[3:0] ? dataArray_15_3_cachedata_MPORT_data : _GEN_6402; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6404 = _GEN_7664 & 4'h4 == EntId[3:0] ? dataArray_15_4_cachedata_MPORT_data : _GEN_6403; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6405 = _GEN_7664 & 4'h5 == EntId[3:0] ? dataArray_15_5_cachedata_MPORT_data : _GEN_6404; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6406 = _GEN_7664 & 4'h6 == EntId[3:0] ? dataArray_15_6_cachedata_MPORT_data : _GEN_6405; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6407 = _GEN_7664 & 4'h7 == EntId[3:0] ? dataArray_15_7_cachedata_MPORT_data : _GEN_6406; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6408 = _GEN_7664 & 4'h8 == EntId[3:0] ? dataArray_15_8_cachedata_MPORT_data : _GEN_6407; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6409 = _GEN_7664 & 4'h9 == EntId[3:0] ? dataArray_15_9_cachedata_MPORT_data : _GEN_6408; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6410 = _GEN_7664 & 4'ha == EntId[3:0] ? dataArray_15_10_cachedata_MPORT_data : _GEN_6409; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6411 = _GEN_7664 & 4'hb == EntId[3:0] ? dataArray_15_11_cachedata_MPORT_data : _GEN_6410; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6412 = _GEN_7664 & 4'hc == EntId[3:0] ? dataArray_15_12_cachedata_MPORT_data : _GEN_6411; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6413 = _GEN_7664 & 4'hd == EntId[3:0] ? dataArray_15_13_cachedata_MPORT_data : _GEN_6412; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6414 = _GEN_7664 & 4'he == EntId[3:0] ? dataArray_15_14_cachedata_MPORT_data : _GEN_6413; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6415 = _GEN_7664 & 4'hf == EntId[3:0] ? dataArray_15_15_cachedata_MPORT_data : _GEN_6414; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6416 = _GEN_7696 & 4'h0 == EntId[3:0] ? dataArray_16_0_cachedata_MPORT_data : _GEN_6415; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6417 = _GEN_7696 & 4'h1 == EntId[3:0] ? dataArray_16_1_cachedata_MPORT_data : _GEN_6416; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6418 = _GEN_7696 & 4'h2 == EntId[3:0] ? dataArray_16_2_cachedata_MPORT_data : _GEN_6417; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6419 = _GEN_7696 & 4'h3 == EntId[3:0] ? dataArray_16_3_cachedata_MPORT_data : _GEN_6418; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6420 = _GEN_7696 & 4'h4 == EntId[3:0] ? dataArray_16_4_cachedata_MPORT_data : _GEN_6419; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6421 = _GEN_7696 & 4'h5 == EntId[3:0] ? dataArray_16_5_cachedata_MPORT_data : _GEN_6420; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6422 = _GEN_7696 & 4'h6 == EntId[3:0] ? dataArray_16_6_cachedata_MPORT_data : _GEN_6421; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6423 = _GEN_7696 & 4'h7 == EntId[3:0] ? dataArray_16_7_cachedata_MPORT_data : _GEN_6422; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6424 = _GEN_7696 & 4'h8 == EntId[3:0] ? dataArray_16_8_cachedata_MPORT_data : _GEN_6423; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6425 = _GEN_7696 & 4'h9 == EntId[3:0] ? dataArray_16_9_cachedata_MPORT_data : _GEN_6424; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6426 = _GEN_7696 & 4'ha == EntId[3:0] ? dataArray_16_10_cachedata_MPORT_data : _GEN_6425; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6427 = _GEN_7696 & 4'hb == EntId[3:0] ? dataArray_16_11_cachedata_MPORT_data : _GEN_6426; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6428 = _GEN_7696 & 4'hc == EntId[3:0] ? dataArray_16_12_cachedata_MPORT_data : _GEN_6427; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6429 = _GEN_7696 & 4'hd == EntId[3:0] ? dataArray_16_13_cachedata_MPORT_data : _GEN_6428; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6430 = _GEN_7696 & 4'he == EntId[3:0] ? dataArray_16_14_cachedata_MPORT_data : _GEN_6429; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6431 = _GEN_7696 & 4'hf == EntId[3:0] ? dataArray_16_15_cachedata_MPORT_data : _GEN_6430; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6432 = _GEN_7728 & 4'h0 == EntId[3:0] ? dataArray_17_0_cachedata_MPORT_data : _GEN_6431; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6433 = _GEN_7728 & 4'h1 == EntId[3:0] ? dataArray_17_1_cachedata_MPORT_data : _GEN_6432; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6434 = _GEN_7728 & 4'h2 == EntId[3:0] ? dataArray_17_2_cachedata_MPORT_data : _GEN_6433; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6435 = _GEN_7728 & 4'h3 == EntId[3:0] ? dataArray_17_3_cachedata_MPORT_data : _GEN_6434; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6436 = _GEN_7728 & 4'h4 == EntId[3:0] ? dataArray_17_4_cachedata_MPORT_data : _GEN_6435; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6437 = _GEN_7728 & 4'h5 == EntId[3:0] ? dataArray_17_5_cachedata_MPORT_data : _GEN_6436; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6438 = _GEN_7728 & 4'h6 == EntId[3:0] ? dataArray_17_6_cachedata_MPORT_data : _GEN_6437; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6439 = _GEN_7728 & 4'h7 == EntId[3:0] ? dataArray_17_7_cachedata_MPORT_data : _GEN_6438; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6440 = _GEN_7728 & 4'h8 == EntId[3:0] ? dataArray_17_8_cachedata_MPORT_data : _GEN_6439; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6441 = _GEN_7728 & 4'h9 == EntId[3:0] ? dataArray_17_9_cachedata_MPORT_data : _GEN_6440; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6442 = _GEN_7728 & 4'ha == EntId[3:0] ? dataArray_17_10_cachedata_MPORT_data : _GEN_6441; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6443 = _GEN_7728 & 4'hb == EntId[3:0] ? dataArray_17_11_cachedata_MPORT_data : _GEN_6442; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6444 = _GEN_7728 & 4'hc == EntId[3:0] ? dataArray_17_12_cachedata_MPORT_data : _GEN_6443; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6445 = _GEN_7728 & 4'hd == EntId[3:0] ? dataArray_17_13_cachedata_MPORT_data : _GEN_6444; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6446 = _GEN_7728 & 4'he == EntId[3:0] ? dataArray_17_14_cachedata_MPORT_data : _GEN_6445; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6447 = _GEN_7728 & 4'hf == EntId[3:0] ? dataArray_17_15_cachedata_MPORT_data : _GEN_6446; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6448 = _GEN_7760 & 4'h0 == EntId[3:0] ? dataArray_18_0_cachedata_MPORT_data : _GEN_6447; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6449 = _GEN_7760 & 4'h1 == EntId[3:0] ? dataArray_18_1_cachedata_MPORT_data : _GEN_6448; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6450 = _GEN_7760 & 4'h2 == EntId[3:0] ? dataArray_18_2_cachedata_MPORT_data : _GEN_6449; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6451 = _GEN_7760 & 4'h3 == EntId[3:0] ? dataArray_18_3_cachedata_MPORT_data : _GEN_6450; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6452 = _GEN_7760 & 4'h4 == EntId[3:0] ? dataArray_18_4_cachedata_MPORT_data : _GEN_6451; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6453 = _GEN_7760 & 4'h5 == EntId[3:0] ? dataArray_18_5_cachedata_MPORT_data : _GEN_6452; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6454 = _GEN_7760 & 4'h6 == EntId[3:0] ? dataArray_18_6_cachedata_MPORT_data : _GEN_6453; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6455 = _GEN_7760 & 4'h7 == EntId[3:0] ? dataArray_18_7_cachedata_MPORT_data : _GEN_6454; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6456 = _GEN_7760 & 4'h8 == EntId[3:0] ? dataArray_18_8_cachedata_MPORT_data : _GEN_6455; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6457 = _GEN_7760 & 4'h9 == EntId[3:0] ? dataArray_18_9_cachedata_MPORT_data : _GEN_6456; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6458 = _GEN_7760 & 4'ha == EntId[3:0] ? dataArray_18_10_cachedata_MPORT_data : _GEN_6457; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6459 = _GEN_7760 & 4'hb == EntId[3:0] ? dataArray_18_11_cachedata_MPORT_data : _GEN_6458; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6460 = _GEN_7760 & 4'hc == EntId[3:0] ? dataArray_18_12_cachedata_MPORT_data : _GEN_6459; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6461 = _GEN_7760 & 4'hd == EntId[3:0] ? dataArray_18_13_cachedata_MPORT_data : _GEN_6460; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6462 = _GEN_7760 & 4'he == EntId[3:0] ? dataArray_18_14_cachedata_MPORT_data : _GEN_6461; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6463 = _GEN_7760 & 4'hf == EntId[3:0] ? dataArray_18_15_cachedata_MPORT_data : _GEN_6462; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6464 = _GEN_7792 & 4'h0 == EntId[3:0] ? dataArray_19_0_cachedata_MPORT_data : _GEN_6463; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6465 = _GEN_7792 & 4'h1 == EntId[3:0] ? dataArray_19_1_cachedata_MPORT_data : _GEN_6464; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6466 = _GEN_7792 & 4'h2 == EntId[3:0] ? dataArray_19_2_cachedata_MPORT_data : _GEN_6465; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6467 = _GEN_7792 & 4'h3 == EntId[3:0] ? dataArray_19_3_cachedata_MPORT_data : _GEN_6466; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6468 = _GEN_7792 & 4'h4 == EntId[3:0] ? dataArray_19_4_cachedata_MPORT_data : _GEN_6467; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6469 = _GEN_7792 & 4'h5 == EntId[3:0] ? dataArray_19_5_cachedata_MPORT_data : _GEN_6468; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6470 = _GEN_7792 & 4'h6 == EntId[3:0] ? dataArray_19_6_cachedata_MPORT_data : _GEN_6469; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6471 = _GEN_7792 & 4'h7 == EntId[3:0] ? dataArray_19_7_cachedata_MPORT_data : _GEN_6470; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6472 = _GEN_7792 & 4'h8 == EntId[3:0] ? dataArray_19_8_cachedata_MPORT_data : _GEN_6471; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6473 = _GEN_7792 & 4'h9 == EntId[3:0] ? dataArray_19_9_cachedata_MPORT_data : _GEN_6472; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6474 = _GEN_7792 & 4'ha == EntId[3:0] ? dataArray_19_10_cachedata_MPORT_data : _GEN_6473; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6475 = _GEN_7792 & 4'hb == EntId[3:0] ? dataArray_19_11_cachedata_MPORT_data : _GEN_6474; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6476 = _GEN_7792 & 4'hc == EntId[3:0] ? dataArray_19_12_cachedata_MPORT_data : _GEN_6475; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6477 = _GEN_7792 & 4'hd == EntId[3:0] ? dataArray_19_13_cachedata_MPORT_data : _GEN_6476; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6478 = _GEN_7792 & 4'he == EntId[3:0] ? dataArray_19_14_cachedata_MPORT_data : _GEN_6477; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6479 = _GEN_7792 & 4'hf == EntId[3:0] ? dataArray_19_15_cachedata_MPORT_data : _GEN_6478; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6480 = _GEN_7824 & 4'h0 == EntId[3:0] ? dataArray_20_0_cachedata_MPORT_data : _GEN_6479; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6481 = _GEN_7824 & 4'h1 == EntId[3:0] ? dataArray_20_1_cachedata_MPORT_data : _GEN_6480; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6482 = _GEN_7824 & 4'h2 == EntId[3:0] ? dataArray_20_2_cachedata_MPORT_data : _GEN_6481; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6483 = _GEN_7824 & 4'h3 == EntId[3:0] ? dataArray_20_3_cachedata_MPORT_data : _GEN_6482; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6484 = _GEN_7824 & 4'h4 == EntId[3:0] ? dataArray_20_4_cachedata_MPORT_data : _GEN_6483; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6485 = _GEN_7824 & 4'h5 == EntId[3:0] ? dataArray_20_5_cachedata_MPORT_data : _GEN_6484; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6486 = _GEN_7824 & 4'h6 == EntId[3:0] ? dataArray_20_6_cachedata_MPORT_data : _GEN_6485; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6487 = _GEN_7824 & 4'h7 == EntId[3:0] ? dataArray_20_7_cachedata_MPORT_data : _GEN_6486; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6488 = _GEN_7824 & 4'h8 == EntId[3:0] ? dataArray_20_8_cachedata_MPORT_data : _GEN_6487; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6489 = _GEN_7824 & 4'h9 == EntId[3:0] ? dataArray_20_9_cachedata_MPORT_data : _GEN_6488; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6490 = _GEN_7824 & 4'ha == EntId[3:0] ? dataArray_20_10_cachedata_MPORT_data : _GEN_6489; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6491 = _GEN_7824 & 4'hb == EntId[3:0] ? dataArray_20_11_cachedata_MPORT_data : _GEN_6490; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6492 = _GEN_7824 & 4'hc == EntId[3:0] ? dataArray_20_12_cachedata_MPORT_data : _GEN_6491; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6493 = _GEN_7824 & 4'hd == EntId[3:0] ? dataArray_20_13_cachedata_MPORT_data : _GEN_6492; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6494 = _GEN_7824 & 4'he == EntId[3:0] ? dataArray_20_14_cachedata_MPORT_data : _GEN_6493; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6495 = _GEN_7824 & 4'hf == EntId[3:0] ? dataArray_20_15_cachedata_MPORT_data : _GEN_6494; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6496 = _GEN_7856 & 4'h0 == EntId[3:0] ? dataArray_21_0_cachedata_MPORT_data : _GEN_6495; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6497 = _GEN_7856 & 4'h1 == EntId[3:0] ? dataArray_21_1_cachedata_MPORT_data : _GEN_6496; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6498 = _GEN_7856 & 4'h2 == EntId[3:0] ? dataArray_21_2_cachedata_MPORT_data : _GEN_6497; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6499 = _GEN_7856 & 4'h3 == EntId[3:0] ? dataArray_21_3_cachedata_MPORT_data : _GEN_6498; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6500 = _GEN_7856 & 4'h4 == EntId[3:0] ? dataArray_21_4_cachedata_MPORT_data : _GEN_6499; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6501 = _GEN_7856 & 4'h5 == EntId[3:0] ? dataArray_21_5_cachedata_MPORT_data : _GEN_6500; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6502 = _GEN_7856 & 4'h6 == EntId[3:0] ? dataArray_21_6_cachedata_MPORT_data : _GEN_6501; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6503 = _GEN_7856 & 4'h7 == EntId[3:0] ? dataArray_21_7_cachedata_MPORT_data : _GEN_6502; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6504 = _GEN_7856 & 4'h8 == EntId[3:0] ? dataArray_21_8_cachedata_MPORT_data : _GEN_6503; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6505 = _GEN_7856 & 4'h9 == EntId[3:0] ? dataArray_21_9_cachedata_MPORT_data : _GEN_6504; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6506 = _GEN_7856 & 4'ha == EntId[3:0] ? dataArray_21_10_cachedata_MPORT_data : _GEN_6505; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6507 = _GEN_7856 & 4'hb == EntId[3:0] ? dataArray_21_11_cachedata_MPORT_data : _GEN_6506; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6508 = _GEN_7856 & 4'hc == EntId[3:0] ? dataArray_21_12_cachedata_MPORT_data : _GEN_6507; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6509 = _GEN_7856 & 4'hd == EntId[3:0] ? dataArray_21_13_cachedata_MPORT_data : _GEN_6508; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6510 = _GEN_7856 & 4'he == EntId[3:0] ? dataArray_21_14_cachedata_MPORT_data : _GEN_6509; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6511 = _GEN_7856 & 4'hf == EntId[3:0] ? dataArray_21_15_cachedata_MPORT_data : _GEN_6510; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6512 = _GEN_7888 & 4'h0 == EntId[3:0] ? dataArray_22_0_cachedata_MPORT_data : _GEN_6511; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6513 = _GEN_7888 & 4'h1 == EntId[3:0] ? dataArray_22_1_cachedata_MPORT_data : _GEN_6512; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6514 = _GEN_7888 & 4'h2 == EntId[3:0] ? dataArray_22_2_cachedata_MPORT_data : _GEN_6513; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6515 = _GEN_7888 & 4'h3 == EntId[3:0] ? dataArray_22_3_cachedata_MPORT_data : _GEN_6514; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6516 = _GEN_7888 & 4'h4 == EntId[3:0] ? dataArray_22_4_cachedata_MPORT_data : _GEN_6515; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6517 = _GEN_7888 & 4'h5 == EntId[3:0] ? dataArray_22_5_cachedata_MPORT_data : _GEN_6516; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6518 = _GEN_7888 & 4'h6 == EntId[3:0] ? dataArray_22_6_cachedata_MPORT_data : _GEN_6517; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6519 = _GEN_7888 & 4'h7 == EntId[3:0] ? dataArray_22_7_cachedata_MPORT_data : _GEN_6518; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6520 = _GEN_7888 & 4'h8 == EntId[3:0] ? dataArray_22_8_cachedata_MPORT_data : _GEN_6519; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6521 = _GEN_7888 & 4'h9 == EntId[3:0] ? dataArray_22_9_cachedata_MPORT_data : _GEN_6520; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6522 = _GEN_7888 & 4'ha == EntId[3:0] ? dataArray_22_10_cachedata_MPORT_data : _GEN_6521; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6523 = _GEN_7888 & 4'hb == EntId[3:0] ? dataArray_22_11_cachedata_MPORT_data : _GEN_6522; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6524 = _GEN_7888 & 4'hc == EntId[3:0] ? dataArray_22_12_cachedata_MPORT_data : _GEN_6523; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6525 = _GEN_7888 & 4'hd == EntId[3:0] ? dataArray_22_13_cachedata_MPORT_data : _GEN_6524; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6526 = _GEN_7888 & 4'he == EntId[3:0] ? dataArray_22_14_cachedata_MPORT_data : _GEN_6525; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6527 = _GEN_7888 & 4'hf == EntId[3:0] ? dataArray_22_15_cachedata_MPORT_data : _GEN_6526; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6528 = _GEN_7920 & 4'h0 == EntId[3:0] ? dataArray_23_0_cachedata_MPORT_data : _GEN_6527; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6529 = _GEN_7920 & 4'h1 == EntId[3:0] ? dataArray_23_1_cachedata_MPORT_data : _GEN_6528; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6530 = _GEN_7920 & 4'h2 == EntId[3:0] ? dataArray_23_2_cachedata_MPORT_data : _GEN_6529; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6531 = _GEN_7920 & 4'h3 == EntId[3:0] ? dataArray_23_3_cachedata_MPORT_data : _GEN_6530; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6532 = _GEN_7920 & 4'h4 == EntId[3:0] ? dataArray_23_4_cachedata_MPORT_data : _GEN_6531; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6533 = _GEN_7920 & 4'h5 == EntId[3:0] ? dataArray_23_5_cachedata_MPORT_data : _GEN_6532; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6534 = _GEN_7920 & 4'h6 == EntId[3:0] ? dataArray_23_6_cachedata_MPORT_data : _GEN_6533; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6535 = _GEN_7920 & 4'h7 == EntId[3:0] ? dataArray_23_7_cachedata_MPORT_data : _GEN_6534; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6536 = _GEN_7920 & 4'h8 == EntId[3:0] ? dataArray_23_8_cachedata_MPORT_data : _GEN_6535; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6537 = _GEN_7920 & 4'h9 == EntId[3:0] ? dataArray_23_9_cachedata_MPORT_data : _GEN_6536; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6538 = _GEN_7920 & 4'ha == EntId[3:0] ? dataArray_23_10_cachedata_MPORT_data : _GEN_6537; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6539 = _GEN_7920 & 4'hb == EntId[3:0] ? dataArray_23_11_cachedata_MPORT_data : _GEN_6538; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6540 = _GEN_7920 & 4'hc == EntId[3:0] ? dataArray_23_12_cachedata_MPORT_data : _GEN_6539; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6541 = _GEN_7920 & 4'hd == EntId[3:0] ? dataArray_23_13_cachedata_MPORT_data : _GEN_6540; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6542 = _GEN_7920 & 4'he == EntId[3:0] ? dataArray_23_14_cachedata_MPORT_data : _GEN_6541; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6543 = _GEN_7920 & 4'hf == EntId[3:0] ? dataArray_23_15_cachedata_MPORT_data : _GEN_6542; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6544 = _GEN_7952 & 4'h0 == EntId[3:0] ? dataArray_24_0_cachedata_MPORT_data : _GEN_6543; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6545 = _GEN_7952 & 4'h1 == EntId[3:0] ? dataArray_24_1_cachedata_MPORT_data : _GEN_6544; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6546 = _GEN_7952 & 4'h2 == EntId[3:0] ? dataArray_24_2_cachedata_MPORT_data : _GEN_6545; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6547 = _GEN_7952 & 4'h3 == EntId[3:0] ? dataArray_24_3_cachedata_MPORT_data : _GEN_6546; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6548 = _GEN_7952 & 4'h4 == EntId[3:0] ? dataArray_24_4_cachedata_MPORT_data : _GEN_6547; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6549 = _GEN_7952 & 4'h5 == EntId[3:0] ? dataArray_24_5_cachedata_MPORT_data : _GEN_6548; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6550 = _GEN_7952 & 4'h6 == EntId[3:0] ? dataArray_24_6_cachedata_MPORT_data : _GEN_6549; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6551 = _GEN_7952 & 4'h7 == EntId[3:0] ? dataArray_24_7_cachedata_MPORT_data : _GEN_6550; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6552 = _GEN_7952 & 4'h8 == EntId[3:0] ? dataArray_24_8_cachedata_MPORT_data : _GEN_6551; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6553 = _GEN_7952 & 4'h9 == EntId[3:0] ? dataArray_24_9_cachedata_MPORT_data : _GEN_6552; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6554 = _GEN_7952 & 4'ha == EntId[3:0] ? dataArray_24_10_cachedata_MPORT_data : _GEN_6553; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6555 = _GEN_7952 & 4'hb == EntId[3:0] ? dataArray_24_11_cachedata_MPORT_data : _GEN_6554; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6556 = _GEN_7952 & 4'hc == EntId[3:0] ? dataArray_24_12_cachedata_MPORT_data : _GEN_6555; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6557 = _GEN_7952 & 4'hd == EntId[3:0] ? dataArray_24_13_cachedata_MPORT_data : _GEN_6556; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6558 = _GEN_7952 & 4'he == EntId[3:0] ? dataArray_24_14_cachedata_MPORT_data : _GEN_6557; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6559 = _GEN_7952 & 4'hf == EntId[3:0] ? dataArray_24_15_cachedata_MPORT_data : _GEN_6558; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6560 = _GEN_7984 & 4'h0 == EntId[3:0] ? dataArray_25_0_cachedata_MPORT_data : _GEN_6559; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6561 = _GEN_7984 & 4'h1 == EntId[3:0] ? dataArray_25_1_cachedata_MPORT_data : _GEN_6560; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6562 = _GEN_7984 & 4'h2 == EntId[3:0] ? dataArray_25_2_cachedata_MPORT_data : _GEN_6561; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6563 = _GEN_7984 & 4'h3 == EntId[3:0] ? dataArray_25_3_cachedata_MPORT_data : _GEN_6562; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6564 = _GEN_7984 & 4'h4 == EntId[3:0] ? dataArray_25_4_cachedata_MPORT_data : _GEN_6563; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6565 = _GEN_7984 & 4'h5 == EntId[3:0] ? dataArray_25_5_cachedata_MPORT_data : _GEN_6564; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6566 = _GEN_7984 & 4'h6 == EntId[3:0] ? dataArray_25_6_cachedata_MPORT_data : _GEN_6565; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6567 = _GEN_7984 & 4'h7 == EntId[3:0] ? dataArray_25_7_cachedata_MPORT_data : _GEN_6566; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6568 = _GEN_7984 & 4'h8 == EntId[3:0] ? dataArray_25_8_cachedata_MPORT_data : _GEN_6567; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6569 = _GEN_7984 & 4'h9 == EntId[3:0] ? dataArray_25_9_cachedata_MPORT_data : _GEN_6568; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6570 = _GEN_7984 & 4'ha == EntId[3:0] ? dataArray_25_10_cachedata_MPORT_data : _GEN_6569; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6571 = _GEN_7984 & 4'hb == EntId[3:0] ? dataArray_25_11_cachedata_MPORT_data : _GEN_6570; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6572 = _GEN_7984 & 4'hc == EntId[3:0] ? dataArray_25_12_cachedata_MPORT_data : _GEN_6571; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6573 = _GEN_7984 & 4'hd == EntId[3:0] ? dataArray_25_13_cachedata_MPORT_data : _GEN_6572; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6574 = _GEN_7984 & 4'he == EntId[3:0] ? dataArray_25_14_cachedata_MPORT_data : _GEN_6573; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6575 = _GEN_7984 & 4'hf == EntId[3:0] ? dataArray_25_15_cachedata_MPORT_data : _GEN_6574; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6576 = _GEN_8016 & 4'h0 == EntId[3:0] ? dataArray_26_0_cachedata_MPORT_data : _GEN_6575; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6577 = _GEN_8016 & 4'h1 == EntId[3:0] ? dataArray_26_1_cachedata_MPORT_data : _GEN_6576; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6578 = _GEN_8016 & 4'h2 == EntId[3:0] ? dataArray_26_2_cachedata_MPORT_data : _GEN_6577; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6579 = _GEN_8016 & 4'h3 == EntId[3:0] ? dataArray_26_3_cachedata_MPORT_data : _GEN_6578; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6580 = _GEN_8016 & 4'h4 == EntId[3:0] ? dataArray_26_4_cachedata_MPORT_data : _GEN_6579; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6581 = _GEN_8016 & 4'h5 == EntId[3:0] ? dataArray_26_5_cachedata_MPORT_data : _GEN_6580; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6582 = _GEN_8016 & 4'h6 == EntId[3:0] ? dataArray_26_6_cachedata_MPORT_data : _GEN_6581; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6583 = _GEN_8016 & 4'h7 == EntId[3:0] ? dataArray_26_7_cachedata_MPORT_data : _GEN_6582; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6584 = _GEN_8016 & 4'h8 == EntId[3:0] ? dataArray_26_8_cachedata_MPORT_data : _GEN_6583; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6585 = _GEN_8016 & 4'h9 == EntId[3:0] ? dataArray_26_9_cachedata_MPORT_data : _GEN_6584; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6586 = _GEN_8016 & 4'ha == EntId[3:0] ? dataArray_26_10_cachedata_MPORT_data : _GEN_6585; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6587 = _GEN_8016 & 4'hb == EntId[3:0] ? dataArray_26_11_cachedata_MPORT_data : _GEN_6586; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6588 = _GEN_8016 & 4'hc == EntId[3:0] ? dataArray_26_12_cachedata_MPORT_data : _GEN_6587; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6589 = _GEN_8016 & 4'hd == EntId[3:0] ? dataArray_26_13_cachedata_MPORT_data : _GEN_6588; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6590 = _GEN_8016 & 4'he == EntId[3:0] ? dataArray_26_14_cachedata_MPORT_data : _GEN_6589; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6591 = _GEN_8016 & 4'hf == EntId[3:0] ? dataArray_26_15_cachedata_MPORT_data : _GEN_6590; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6592 = _GEN_8048 & 4'h0 == EntId[3:0] ? dataArray_27_0_cachedata_MPORT_data : _GEN_6591; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6593 = _GEN_8048 & 4'h1 == EntId[3:0] ? dataArray_27_1_cachedata_MPORT_data : _GEN_6592; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6594 = _GEN_8048 & 4'h2 == EntId[3:0] ? dataArray_27_2_cachedata_MPORT_data : _GEN_6593; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6595 = _GEN_8048 & 4'h3 == EntId[3:0] ? dataArray_27_3_cachedata_MPORT_data : _GEN_6594; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6596 = _GEN_8048 & 4'h4 == EntId[3:0] ? dataArray_27_4_cachedata_MPORT_data : _GEN_6595; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6597 = _GEN_8048 & 4'h5 == EntId[3:0] ? dataArray_27_5_cachedata_MPORT_data : _GEN_6596; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6598 = _GEN_8048 & 4'h6 == EntId[3:0] ? dataArray_27_6_cachedata_MPORT_data : _GEN_6597; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6599 = _GEN_8048 & 4'h7 == EntId[3:0] ? dataArray_27_7_cachedata_MPORT_data : _GEN_6598; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6600 = _GEN_8048 & 4'h8 == EntId[3:0] ? dataArray_27_8_cachedata_MPORT_data : _GEN_6599; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6601 = _GEN_8048 & 4'h9 == EntId[3:0] ? dataArray_27_9_cachedata_MPORT_data : _GEN_6600; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6602 = _GEN_8048 & 4'ha == EntId[3:0] ? dataArray_27_10_cachedata_MPORT_data : _GEN_6601; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6603 = _GEN_8048 & 4'hb == EntId[3:0] ? dataArray_27_11_cachedata_MPORT_data : _GEN_6602; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6604 = _GEN_8048 & 4'hc == EntId[3:0] ? dataArray_27_12_cachedata_MPORT_data : _GEN_6603; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6605 = _GEN_8048 & 4'hd == EntId[3:0] ? dataArray_27_13_cachedata_MPORT_data : _GEN_6604; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6606 = _GEN_8048 & 4'he == EntId[3:0] ? dataArray_27_14_cachedata_MPORT_data : _GEN_6605; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6607 = _GEN_8048 & 4'hf == EntId[3:0] ? dataArray_27_15_cachedata_MPORT_data : _GEN_6606; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6608 = _GEN_8080 & 4'h0 == EntId[3:0] ? dataArray_28_0_cachedata_MPORT_data : _GEN_6607; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6609 = _GEN_8080 & 4'h1 == EntId[3:0] ? dataArray_28_1_cachedata_MPORT_data : _GEN_6608; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6610 = _GEN_8080 & 4'h2 == EntId[3:0] ? dataArray_28_2_cachedata_MPORT_data : _GEN_6609; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6611 = _GEN_8080 & 4'h3 == EntId[3:0] ? dataArray_28_3_cachedata_MPORT_data : _GEN_6610; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6612 = _GEN_8080 & 4'h4 == EntId[3:0] ? dataArray_28_4_cachedata_MPORT_data : _GEN_6611; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6613 = _GEN_8080 & 4'h5 == EntId[3:0] ? dataArray_28_5_cachedata_MPORT_data : _GEN_6612; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6614 = _GEN_8080 & 4'h6 == EntId[3:0] ? dataArray_28_6_cachedata_MPORT_data : _GEN_6613; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6615 = _GEN_8080 & 4'h7 == EntId[3:0] ? dataArray_28_7_cachedata_MPORT_data : _GEN_6614; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6616 = _GEN_8080 & 4'h8 == EntId[3:0] ? dataArray_28_8_cachedata_MPORT_data : _GEN_6615; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6617 = _GEN_8080 & 4'h9 == EntId[3:0] ? dataArray_28_9_cachedata_MPORT_data : _GEN_6616; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6618 = _GEN_8080 & 4'ha == EntId[3:0] ? dataArray_28_10_cachedata_MPORT_data : _GEN_6617; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6619 = _GEN_8080 & 4'hb == EntId[3:0] ? dataArray_28_11_cachedata_MPORT_data : _GEN_6618; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6620 = _GEN_8080 & 4'hc == EntId[3:0] ? dataArray_28_12_cachedata_MPORT_data : _GEN_6619; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6621 = _GEN_8080 & 4'hd == EntId[3:0] ? dataArray_28_13_cachedata_MPORT_data : _GEN_6620; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6622 = _GEN_8080 & 4'he == EntId[3:0] ? dataArray_28_14_cachedata_MPORT_data : _GEN_6621; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6623 = _GEN_8080 & 4'hf == EntId[3:0] ? dataArray_28_15_cachedata_MPORT_data : _GEN_6622; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6624 = _GEN_8112 & 4'h0 == EntId[3:0] ? dataArray_29_0_cachedata_MPORT_data : _GEN_6623; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6625 = _GEN_8112 & 4'h1 == EntId[3:0] ? dataArray_29_1_cachedata_MPORT_data : _GEN_6624; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6626 = _GEN_8112 & 4'h2 == EntId[3:0] ? dataArray_29_2_cachedata_MPORT_data : _GEN_6625; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6627 = _GEN_8112 & 4'h3 == EntId[3:0] ? dataArray_29_3_cachedata_MPORT_data : _GEN_6626; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6628 = _GEN_8112 & 4'h4 == EntId[3:0] ? dataArray_29_4_cachedata_MPORT_data : _GEN_6627; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6629 = _GEN_8112 & 4'h5 == EntId[3:0] ? dataArray_29_5_cachedata_MPORT_data : _GEN_6628; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6630 = _GEN_8112 & 4'h6 == EntId[3:0] ? dataArray_29_6_cachedata_MPORT_data : _GEN_6629; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6631 = _GEN_8112 & 4'h7 == EntId[3:0] ? dataArray_29_7_cachedata_MPORT_data : _GEN_6630; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6632 = _GEN_8112 & 4'h8 == EntId[3:0] ? dataArray_29_8_cachedata_MPORT_data : _GEN_6631; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6633 = _GEN_8112 & 4'h9 == EntId[3:0] ? dataArray_29_9_cachedata_MPORT_data : _GEN_6632; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6634 = _GEN_8112 & 4'ha == EntId[3:0] ? dataArray_29_10_cachedata_MPORT_data : _GEN_6633; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6635 = _GEN_8112 & 4'hb == EntId[3:0] ? dataArray_29_11_cachedata_MPORT_data : _GEN_6634; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6636 = _GEN_8112 & 4'hc == EntId[3:0] ? dataArray_29_12_cachedata_MPORT_data : _GEN_6635; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6637 = _GEN_8112 & 4'hd == EntId[3:0] ? dataArray_29_13_cachedata_MPORT_data : _GEN_6636; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6638 = _GEN_8112 & 4'he == EntId[3:0] ? dataArray_29_14_cachedata_MPORT_data : _GEN_6637; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6639 = _GEN_8112 & 4'hf == EntId[3:0] ? dataArray_29_15_cachedata_MPORT_data : _GEN_6638; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6640 = _GEN_8144 & 4'h0 == EntId[3:0] ? dataArray_30_0_cachedata_MPORT_data : _GEN_6639; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6641 = _GEN_8144 & 4'h1 == EntId[3:0] ? dataArray_30_1_cachedata_MPORT_data : _GEN_6640; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6642 = _GEN_8144 & 4'h2 == EntId[3:0] ? dataArray_30_2_cachedata_MPORT_data : _GEN_6641; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6643 = _GEN_8144 & 4'h3 == EntId[3:0] ? dataArray_30_3_cachedata_MPORT_data : _GEN_6642; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6644 = _GEN_8144 & 4'h4 == EntId[3:0] ? dataArray_30_4_cachedata_MPORT_data : _GEN_6643; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6645 = _GEN_8144 & 4'h5 == EntId[3:0] ? dataArray_30_5_cachedata_MPORT_data : _GEN_6644; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6646 = _GEN_8144 & 4'h6 == EntId[3:0] ? dataArray_30_6_cachedata_MPORT_data : _GEN_6645; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6647 = _GEN_8144 & 4'h7 == EntId[3:0] ? dataArray_30_7_cachedata_MPORT_data : _GEN_6646; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6648 = _GEN_8144 & 4'h8 == EntId[3:0] ? dataArray_30_8_cachedata_MPORT_data : _GEN_6647; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6649 = _GEN_8144 & 4'h9 == EntId[3:0] ? dataArray_30_9_cachedata_MPORT_data : _GEN_6648; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6650 = _GEN_8144 & 4'ha == EntId[3:0] ? dataArray_30_10_cachedata_MPORT_data : _GEN_6649; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6651 = _GEN_8144 & 4'hb == EntId[3:0] ? dataArray_30_11_cachedata_MPORT_data : _GEN_6650; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6652 = _GEN_8144 & 4'hc == EntId[3:0] ? dataArray_30_12_cachedata_MPORT_data : _GEN_6651; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6653 = _GEN_8144 & 4'hd == EntId[3:0] ? dataArray_30_13_cachedata_MPORT_data : _GEN_6652; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6654 = _GEN_8144 & 4'he == EntId[3:0] ? dataArray_30_14_cachedata_MPORT_data : _GEN_6653; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6655 = _GEN_8144 & 4'hf == EntId[3:0] ? dataArray_30_15_cachedata_MPORT_data : _GEN_6654; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6656 = _GEN_8176 & 4'h0 == EntId[3:0] ? dataArray_31_0_cachedata_MPORT_data : _GEN_6655; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6657 = _GEN_8176 & 4'h1 == EntId[3:0] ? dataArray_31_1_cachedata_MPORT_data : _GEN_6656; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6658 = _GEN_8176 & 4'h2 == EntId[3:0] ? dataArray_31_2_cachedata_MPORT_data : _GEN_6657; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6659 = _GEN_8176 & 4'h3 == EntId[3:0] ? dataArray_31_3_cachedata_MPORT_data : _GEN_6658; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6660 = _GEN_8176 & 4'h4 == EntId[3:0] ? dataArray_31_4_cachedata_MPORT_data : _GEN_6659; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6661 = _GEN_8176 & 4'h5 == EntId[3:0] ? dataArray_31_5_cachedata_MPORT_data : _GEN_6660; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6662 = _GEN_8176 & 4'h6 == EntId[3:0] ? dataArray_31_6_cachedata_MPORT_data : _GEN_6661; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6663 = _GEN_8176 & 4'h7 == EntId[3:0] ? dataArray_31_7_cachedata_MPORT_data : _GEN_6662; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6664 = _GEN_8176 & 4'h8 == EntId[3:0] ? dataArray_31_8_cachedata_MPORT_data : _GEN_6663; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6665 = _GEN_8176 & 4'h9 == EntId[3:0] ? dataArray_31_9_cachedata_MPORT_data : _GEN_6664; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6666 = _GEN_8176 & 4'ha == EntId[3:0] ? dataArray_31_10_cachedata_MPORT_data : _GEN_6665; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6667 = _GEN_8176 & 4'hb == EntId[3:0] ? dataArray_31_11_cachedata_MPORT_data : _GEN_6666; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6668 = _GEN_8176 & 4'hc == EntId[3:0] ? dataArray_31_12_cachedata_MPORT_data : _GEN_6667; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6669 = _GEN_8176 & 4'hd == EntId[3:0] ? dataArray_31_13_cachedata_MPORT_data : _GEN_6668; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6670 = _GEN_8176 & 4'he == EntId[3:0] ? dataArray_31_14_cachedata_MPORT_data : _GEN_6669; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6671 = _GEN_8176 & 4'hf == EntId[3:0] ? dataArray_31_15_cachedata_MPORT_data : _GEN_6670; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6672 = _GEN_8208 & 4'h0 == EntId[3:0] ? dataArray_32_0_cachedata_MPORT_data : _GEN_6671; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6673 = _GEN_8208 & 4'h1 == EntId[3:0] ? dataArray_32_1_cachedata_MPORT_data : _GEN_6672; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6674 = _GEN_8208 & 4'h2 == EntId[3:0] ? dataArray_32_2_cachedata_MPORT_data : _GEN_6673; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6675 = _GEN_8208 & 4'h3 == EntId[3:0] ? dataArray_32_3_cachedata_MPORT_data : _GEN_6674; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6676 = _GEN_8208 & 4'h4 == EntId[3:0] ? dataArray_32_4_cachedata_MPORT_data : _GEN_6675; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6677 = _GEN_8208 & 4'h5 == EntId[3:0] ? dataArray_32_5_cachedata_MPORT_data : _GEN_6676; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6678 = _GEN_8208 & 4'h6 == EntId[3:0] ? dataArray_32_6_cachedata_MPORT_data : _GEN_6677; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6679 = _GEN_8208 & 4'h7 == EntId[3:0] ? dataArray_32_7_cachedata_MPORT_data : _GEN_6678; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6680 = _GEN_8208 & 4'h8 == EntId[3:0] ? dataArray_32_8_cachedata_MPORT_data : _GEN_6679; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6681 = _GEN_8208 & 4'h9 == EntId[3:0] ? dataArray_32_9_cachedata_MPORT_data : _GEN_6680; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6682 = _GEN_8208 & 4'ha == EntId[3:0] ? dataArray_32_10_cachedata_MPORT_data : _GEN_6681; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6683 = _GEN_8208 & 4'hb == EntId[3:0] ? dataArray_32_11_cachedata_MPORT_data : _GEN_6682; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6684 = _GEN_8208 & 4'hc == EntId[3:0] ? dataArray_32_12_cachedata_MPORT_data : _GEN_6683; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6685 = _GEN_8208 & 4'hd == EntId[3:0] ? dataArray_32_13_cachedata_MPORT_data : _GEN_6684; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6686 = _GEN_8208 & 4'he == EntId[3:0] ? dataArray_32_14_cachedata_MPORT_data : _GEN_6685; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6687 = _GEN_8208 & 4'hf == EntId[3:0] ? dataArray_32_15_cachedata_MPORT_data : _GEN_6686; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6688 = _GEN_8240 & 4'h0 == EntId[3:0] ? dataArray_33_0_cachedata_MPORT_data : _GEN_6687; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6689 = _GEN_8240 & 4'h1 == EntId[3:0] ? dataArray_33_1_cachedata_MPORT_data : _GEN_6688; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6690 = _GEN_8240 & 4'h2 == EntId[3:0] ? dataArray_33_2_cachedata_MPORT_data : _GEN_6689; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6691 = _GEN_8240 & 4'h3 == EntId[3:0] ? dataArray_33_3_cachedata_MPORT_data : _GEN_6690; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6692 = _GEN_8240 & 4'h4 == EntId[3:0] ? dataArray_33_4_cachedata_MPORT_data : _GEN_6691; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6693 = _GEN_8240 & 4'h5 == EntId[3:0] ? dataArray_33_5_cachedata_MPORT_data : _GEN_6692; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6694 = _GEN_8240 & 4'h6 == EntId[3:0] ? dataArray_33_6_cachedata_MPORT_data : _GEN_6693; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6695 = _GEN_8240 & 4'h7 == EntId[3:0] ? dataArray_33_7_cachedata_MPORT_data : _GEN_6694; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6696 = _GEN_8240 & 4'h8 == EntId[3:0] ? dataArray_33_8_cachedata_MPORT_data : _GEN_6695; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6697 = _GEN_8240 & 4'h9 == EntId[3:0] ? dataArray_33_9_cachedata_MPORT_data : _GEN_6696; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6698 = _GEN_8240 & 4'ha == EntId[3:0] ? dataArray_33_10_cachedata_MPORT_data : _GEN_6697; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6699 = _GEN_8240 & 4'hb == EntId[3:0] ? dataArray_33_11_cachedata_MPORT_data : _GEN_6698; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6700 = _GEN_8240 & 4'hc == EntId[3:0] ? dataArray_33_12_cachedata_MPORT_data : _GEN_6699; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6701 = _GEN_8240 & 4'hd == EntId[3:0] ? dataArray_33_13_cachedata_MPORT_data : _GEN_6700; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6702 = _GEN_8240 & 4'he == EntId[3:0] ? dataArray_33_14_cachedata_MPORT_data : _GEN_6701; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6703 = _GEN_8240 & 4'hf == EntId[3:0] ? dataArray_33_15_cachedata_MPORT_data : _GEN_6702; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6704 = _GEN_8272 & 4'h0 == EntId[3:0] ? dataArray_34_0_cachedata_MPORT_data : _GEN_6703; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6705 = _GEN_8272 & 4'h1 == EntId[3:0] ? dataArray_34_1_cachedata_MPORT_data : _GEN_6704; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6706 = _GEN_8272 & 4'h2 == EntId[3:0] ? dataArray_34_2_cachedata_MPORT_data : _GEN_6705; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6707 = _GEN_8272 & 4'h3 == EntId[3:0] ? dataArray_34_3_cachedata_MPORT_data : _GEN_6706; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6708 = _GEN_8272 & 4'h4 == EntId[3:0] ? dataArray_34_4_cachedata_MPORT_data : _GEN_6707; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6709 = _GEN_8272 & 4'h5 == EntId[3:0] ? dataArray_34_5_cachedata_MPORT_data : _GEN_6708; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6710 = _GEN_8272 & 4'h6 == EntId[3:0] ? dataArray_34_6_cachedata_MPORT_data : _GEN_6709; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6711 = _GEN_8272 & 4'h7 == EntId[3:0] ? dataArray_34_7_cachedata_MPORT_data : _GEN_6710; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6712 = _GEN_8272 & 4'h8 == EntId[3:0] ? dataArray_34_8_cachedata_MPORT_data : _GEN_6711; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6713 = _GEN_8272 & 4'h9 == EntId[3:0] ? dataArray_34_9_cachedata_MPORT_data : _GEN_6712; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6714 = _GEN_8272 & 4'ha == EntId[3:0] ? dataArray_34_10_cachedata_MPORT_data : _GEN_6713; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6715 = _GEN_8272 & 4'hb == EntId[3:0] ? dataArray_34_11_cachedata_MPORT_data : _GEN_6714; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6716 = _GEN_8272 & 4'hc == EntId[3:0] ? dataArray_34_12_cachedata_MPORT_data : _GEN_6715; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6717 = _GEN_8272 & 4'hd == EntId[3:0] ? dataArray_34_13_cachedata_MPORT_data : _GEN_6716; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6718 = _GEN_8272 & 4'he == EntId[3:0] ? dataArray_34_14_cachedata_MPORT_data : _GEN_6717; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6719 = _GEN_8272 & 4'hf == EntId[3:0] ? dataArray_34_15_cachedata_MPORT_data : _GEN_6718; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6720 = _GEN_8304 & 4'h0 == EntId[3:0] ? dataArray_35_0_cachedata_MPORT_data : _GEN_6719; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6721 = _GEN_8304 & 4'h1 == EntId[3:0] ? dataArray_35_1_cachedata_MPORT_data : _GEN_6720; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6722 = _GEN_8304 & 4'h2 == EntId[3:0] ? dataArray_35_2_cachedata_MPORT_data : _GEN_6721; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6723 = _GEN_8304 & 4'h3 == EntId[3:0] ? dataArray_35_3_cachedata_MPORT_data : _GEN_6722; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6724 = _GEN_8304 & 4'h4 == EntId[3:0] ? dataArray_35_4_cachedata_MPORT_data : _GEN_6723; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6725 = _GEN_8304 & 4'h5 == EntId[3:0] ? dataArray_35_5_cachedata_MPORT_data : _GEN_6724; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6726 = _GEN_8304 & 4'h6 == EntId[3:0] ? dataArray_35_6_cachedata_MPORT_data : _GEN_6725; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6727 = _GEN_8304 & 4'h7 == EntId[3:0] ? dataArray_35_7_cachedata_MPORT_data : _GEN_6726; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6728 = _GEN_8304 & 4'h8 == EntId[3:0] ? dataArray_35_8_cachedata_MPORT_data : _GEN_6727; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6729 = _GEN_8304 & 4'h9 == EntId[3:0] ? dataArray_35_9_cachedata_MPORT_data : _GEN_6728; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6730 = _GEN_8304 & 4'ha == EntId[3:0] ? dataArray_35_10_cachedata_MPORT_data : _GEN_6729; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6731 = _GEN_8304 & 4'hb == EntId[3:0] ? dataArray_35_11_cachedata_MPORT_data : _GEN_6730; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6732 = _GEN_8304 & 4'hc == EntId[3:0] ? dataArray_35_12_cachedata_MPORT_data : _GEN_6731; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6733 = _GEN_8304 & 4'hd == EntId[3:0] ? dataArray_35_13_cachedata_MPORT_data : _GEN_6732; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6734 = _GEN_8304 & 4'he == EntId[3:0] ? dataArray_35_14_cachedata_MPORT_data : _GEN_6733; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6735 = _GEN_8304 & 4'hf == EntId[3:0] ? dataArray_35_15_cachedata_MPORT_data : _GEN_6734; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6736 = _GEN_8336 & 4'h0 == EntId[3:0] ? dataArray_36_0_cachedata_MPORT_data : _GEN_6735; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6737 = _GEN_8336 & 4'h1 == EntId[3:0] ? dataArray_36_1_cachedata_MPORT_data : _GEN_6736; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6738 = _GEN_8336 & 4'h2 == EntId[3:0] ? dataArray_36_2_cachedata_MPORT_data : _GEN_6737; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6739 = _GEN_8336 & 4'h3 == EntId[3:0] ? dataArray_36_3_cachedata_MPORT_data : _GEN_6738; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6740 = _GEN_8336 & 4'h4 == EntId[3:0] ? dataArray_36_4_cachedata_MPORT_data : _GEN_6739; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6741 = _GEN_8336 & 4'h5 == EntId[3:0] ? dataArray_36_5_cachedata_MPORT_data : _GEN_6740; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6742 = _GEN_8336 & 4'h6 == EntId[3:0] ? dataArray_36_6_cachedata_MPORT_data : _GEN_6741; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6743 = _GEN_8336 & 4'h7 == EntId[3:0] ? dataArray_36_7_cachedata_MPORT_data : _GEN_6742; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6744 = _GEN_8336 & 4'h8 == EntId[3:0] ? dataArray_36_8_cachedata_MPORT_data : _GEN_6743; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6745 = _GEN_8336 & 4'h9 == EntId[3:0] ? dataArray_36_9_cachedata_MPORT_data : _GEN_6744; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6746 = _GEN_8336 & 4'ha == EntId[3:0] ? dataArray_36_10_cachedata_MPORT_data : _GEN_6745; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6747 = _GEN_8336 & 4'hb == EntId[3:0] ? dataArray_36_11_cachedata_MPORT_data : _GEN_6746; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6748 = _GEN_8336 & 4'hc == EntId[3:0] ? dataArray_36_12_cachedata_MPORT_data : _GEN_6747; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6749 = _GEN_8336 & 4'hd == EntId[3:0] ? dataArray_36_13_cachedata_MPORT_data : _GEN_6748; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6750 = _GEN_8336 & 4'he == EntId[3:0] ? dataArray_36_14_cachedata_MPORT_data : _GEN_6749; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6751 = _GEN_8336 & 4'hf == EntId[3:0] ? dataArray_36_15_cachedata_MPORT_data : _GEN_6750; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6752 = _GEN_8368 & 4'h0 == EntId[3:0] ? dataArray_37_0_cachedata_MPORT_data : _GEN_6751; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6753 = _GEN_8368 & 4'h1 == EntId[3:0] ? dataArray_37_1_cachedata_MPORT_data : _GEN_6752; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6754 = _GEN_8368 & 4'h2 == EntId[3:0] ? dataArray_37_2_cachedata_MPORT_data : _GEN_6753; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6755 = _GEN_8368 & 4'h3 == EntId[3:0] ? dataArray_37_3_cachedata_MPORT_data : _GEN_6754; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6756 = _GEN_8368 & 4'h4 == EntId[3:0] ? dataArray_37_4_cachedata_MPORT_data : _GEN_6755; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6757 = _GEN_8368 & 4'h5 == EntId[3:0] ? dataArray_37_5_cachedata_MPORT_data : _GEN_6756; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6758 = _GEN_8368 & 4'h6 == EntId[3:0] ? dataArray_37_6_cachedata_MPORT_data : _GEN_6757; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6759 = _GEN_8368 & 4'h7 == EntId[3:0] ? dataArray_37_7_cachedata_MPORT_data : _GEN_6758; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6760 = _GEN_8368 & 4'h8 == EntId[3:0] ? dataArray_37_8_cachedata_MPORT_data : _GEN_6759; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6761 = _GEN_8368 & 4'h9 == EntId[3:0] ? dataArray_37_9_cachedata_MPORT_data : _GEN_6760; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6762 = _GEN_8368 & 4'ha == EntId[3:0] ? dataArray_37_10_cachedata_MPORT_data : _GEN_6761; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6763 = _GEN_8368 & 4'hb == EntId[3:0] ? dataArray_37_11_cachedata_MPORT_data : _GEN_6762; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6764 = _GEN_8368 & 4'hc == EntId[3:0] ? dataArray_37_12_cachedata_MPORT_data : _GEN_6763; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6765 = _GEN_8368 & 4'hd == EntId[3:0] ? dataArray_37_13_cachedata_MPORT_data : _GEN_6764; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6766 = _GEN_8368 & 4'he == EntId[3:0] ? dataArray_37_14_cachedata_MPORT_data : _GEN_6765; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6767 = _GEN_8368 & 4'hf == EntId[3:0] ? dataArray_37_15_cachedata_MPORT_data : _GEN_6766; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6768 = _GEN_8400 & 4'h0 == EntId[3:0] ? dataArray_38_0_cachedata_MPORT_data : _GEN_6767; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6769 = _GEN_8400 & 4'h1 == EntId[3:0] ? dataArray_38_1_cachedata_MPORT_data : _GEN_6768; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6770 = _GEN_8400 & 4'h2 == EntId[3:0] ? dataArray_38_2_cachedata_MPORT_data : _GEN_6769; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6771 = _GEN_8400 & 4'h3 == EntId[3:0] ? dataArray_38_3_cachedata_MPORT_data : _GEN_6770; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6772 = _GEN_8400 & 4'h4 == EntId[3:0] ? dataArray_38_4_cachedata_MPORT_data : _GEN_6771; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6773 = _GEN_8400 & 4'h5 == EntId[3:0] ? dataArray_38_5_cachedata_MPORT_data : _GEN_6772; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6774 = _GEN_8400 & 4'h6 == EntId[3:0] ? dataArray_38_6_cachedata_MPORT_data : _GEN_6773; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6775 = _GEN_8400 & 4'h7 == EntId[3:0] ? dataArray_38_7_cachedata_MPORT_data : _GEN_6774; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6776 = _GEN_8400 & 4'h8 == EntId[3:0] ? dataArray_38_8_cachedata_MPORT_data : _GEN_6775; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6777 = _GEN_8400 & 4'h9 == EntId[3:0] ? dataArray_38_9_cachedata_MPORT_data : _GEN_6776; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6778 = _GEN_8400 & 4'ha == EntId[3:0] ? dataArray_38_10_cachedata_MPORT_data : _GEN_6777; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6779 = _GEN_8400 & 4'hb == EntId[3:0] ? dataArray_38_11_cachedata_MPORT_data : _GEN_6778; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6780 = _GEN_8400 & 4'hc == EntId[3:0] ? dataArray_38_12_cachedata_MPORT_data : _GEN_6779; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6781 = _GEN_8400 & 4'hd == EntId[3:0] ? dataArray_38_13_cachedata_MPORT_data : _GEN_6780; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6782 = _GEN_8400 & 4'he == EntId[3:0] ? dataArray_38_14_cachedata_MPORT_data : _GEN_6781; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6783 = _GEN_8400 & 4'hf == EntId[3:0] ? dataArray_38_15_cachedata_MPORT_data : _GEN_6782; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6784 = _GEN_8432 & 4'h0 == EntId[3:0] ? dataArray_39_0_cachedata_MPORT_data : _GEN_6783; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6785 = _GEN_8432 & 4'h1 == EntId[3:0] ? dataArray_39_1_cachedata_MPORT_data : _GEN_6784; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6786 = _GEN_8432 & 4'h2 == EntId[3:0] ? dataArray_39_2_cachedata_MPORT_data : _GEN_6785; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6787 = _GEN_8432 & 4'h3 == EntId[3:0] ? dataArray_39_3_cachedata_MPORT_data : _GEN_6786; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6788 = _GEN_8432 & 4'h4 == EntId[3:0] ? dataArray_39_4_cachedata_MPORT_data : _GEN_6787; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6789 = _GEN_8432 & 4'h5 == EntId[3:0] ? dataArray_39_5_cachedata_MPORT_data : _GEN_6788; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6790 = _GEN_8432 & 4'h6 == EntId[3:0] ? dataArray_39_6_cachedata_MPORT_data : _GEN_6789; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6791 = _GEN_8432 & 4'h7 == EntId[3:0] ? dataArray_39_7_cachedata_MPORT_data : _GEN_6790; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6792 = _GEN_8432 & 4'h8 == EntId[3:0] ? dataArray_39_8_cachedata_MPORT_data : _GEN_6791; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6793 = _GEN_8432 & 4'h9 == EntId[3:0] ? dataArray_39_9_cachedata_MPORT_data : _GEN_6792; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6794 = _GEN_8432 & 4'ha == EntId[3:0] ? dataArray_39_10_cachedata_MPORT_data : _GEN_6793; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6795 = _GEN_8432 & 4'hb == EntId[3:0] ? dataArray_39_11_cachedata_MPORT_data : _GEN_6794; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6796 = _GEN_8432 & 4'hc == EntId[3:0] ? dataArray_39_12_cachedata_MPORT_data : _GEN_6795; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6797 = _GEN_8432 & 4'hd == EntId[3:0] ? dataArray_39_13_cachedata_MPORT_data : _GEN_6796; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6798 = _GEN_8432 & 4'he == EntId[3:0] ? dataArray_39_14_cachedata_MPORT_data : _GEN_6797; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6799 = _GEN_8432 & 4'hf == EntId[3:0] ? dataArray_39_15_cachedata_MPORT_data : _GEN_6798; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6800 = _GEN_8464 & 4'h0 == EntId[3:0] ? dataArray_40_0_cachedata_MPORT_data : _GEN_6799; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6801 = _GEN_8464 & 4'h1 == EntId[3:0] ? dataArray_40_1_cachedata_MPORT_data : _GEN_6800; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6802 = _GEN_8464 & 4'h2 == EntId[3:0] ? dataArray_40_2_cachedata_MPORT_data : _GEN_6801; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6803 = _GEN_8464 & 4'h3 == EntId[3:0] ? dataArray_40_3_cachedata_MPORT_data : _GEN_6802; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6804 = _GEN_8464 & 4'h4 == EntId[3:0] ? dataArray_40_4_cachedata_MPORT_data : _GEN_6803; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6805 = _GEN_8464 & 4'h5 == EntId[3:0] ? dataArray_40_5_cachedata_MPORT_data : _GEN_6804; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6806 = _GEN_8464 & 4'h6 == EntId[3:0] ? dataArray_40_6_cachedata_MPORT_data : _GEN_6805; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6807 = _GEN_8464 & 4'h7 == EntId[3:0] ? dataArray_40_7_cachedata_MPORT_data : _GEN_6806; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6808 = _GEN_8464 & 4'h8 == EntId[3:0] ? dataArray_40_8_cachedata_MPORT_data : _GEN_6807; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6809 = _GEN_8464 & 4'h9 == EntId[3:0] ? dataArray_40_9_cachedata_MPORT_data : _GEN_6808; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6810 = _GEN_8464 & 4'ha == EntId[3:0] ? dataArray_40_10_cachedata_MPORT_data : _GEN_6809; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6811 = _GEN_8464 & 4'hb == EntId[3:0] ? dataArray_40_11_cachedata_MPORT_data : _GEN_6810; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6812 = _GEN_8464 & 4'hc == EntId[3:0] ? dataArray_40_12_cachedata_MPORT_data : _GEN_6811; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6813 = _GEN_8464 & 4'hd == EntId[3:0] ? dataArray_40_13_cachedata_MPORT_data : _GEN_6812; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6814 = _GEN_8464 & 4'he == EntId[3:0] ? dataArray_40_14_cachedata_MPORT_data : _GEN_6813; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6815 = _GEN_8464 & 4'hf == EntId[3:0] ? dataArray_40_15_cachedata_MPORT_data : _GEN_6814; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6816 = _GEN_8496 & 4'h0 == EntId[3:0] ? dataArray_41_0_cachedata_MPORT_data : _GEN_6815; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6817 = _GEN_8496 & 4'h1 == EntId[3:0] ? dataArray_41_1_cachedata_MPORT_data : _GEN_6816; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6818 = _GEN_8496 & 4'h2 == EntId[3:0] ? dataArray_41_2_cachedata_MPORT_data : _GEN_6817; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6819 = _GEN_8496 & 4'h3 == EntId[3:0] ? dataArray_41_3_cachedata_MPORT_data : _GEN_6818; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6820 = _GEN_8496 & 4'h4 == EntId[3:0] ? dataArray_41_4_cachedata_MPORT_data : _GEN_6819; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6821 = _GEN_8496 & 4'h5 == EntId[3:0] ? dataArray_41_5_cachedata_MPORT_data : _GEN_6820; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6822 = _GEN_8496 & 4'h6 == EntId[3:0] ? dataArray_41_6_cachedata_MPORT_data : _GEN_6821; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6823 = _GEN_8496 & 4'h7 == EntId[3:0] ? dataArray_41_7_cachedata_MPORT_data : _GEN_6822; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6824 = _GEN_8496 & 4'h8 == EntId[3:0] ? dataArray_41_8_cachedata_MPORT_data : _GEN_6823; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6825 = _GEN_8496 & 4'h9 == EntId[3:0] ? dataArray_41_9_cachedata_MPORT_data : _GEN_6824; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6826 = _GEN_8496 & 4'ha == EntId[3:0] ? dataArray_41_10_cachedata_MPORT_data : _GEN_6825; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6827 = _GEN_8496 & 4'hb == EntId[3:0] ? dataArray_41_11_cachedata_MPORT_data : _GEN_6826; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6828 = _GEN_8496 & 4'hc == EntId[3:0] ? dataArray_41_12_cachedata_MPORT_data : _GEN_6827; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6829 = _GEN_8496 & 4'hd == EntId[3:0] ? dataArray_41_13_cachedata_MPORT_data : _GEN_6828; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6830 = _GEN_8496 & 4'he == EntId[3:0] ? dataArray_41_14_cachedata_MPORT_data : _GEN_6829; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6831 = _GEN_8496 & 4'hf == EntId[3:0] ? dataArray_41_15_cachedata_MPORT_data : _GEN_6830; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6832 = _GEN_8528 & 4'h0 == EntId[3:0] ? dataArray_42_0_cachedata_MPORT_data : _GEN_6831; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6833 = _GEN_8528 & 4'h1 == EntId[3:0] ? dataArray_42_1_cachedata_MPORT_data : _GEN_6832; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6834 = _GEN_8528 & 4'h2 == EntId[3:0] ? dataArray_42_2_cachedata_MPORT_data : _GEN_6833; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6835 = _GEN_8528 & 4'h3 == EntId[3:0] ? dataArray_42_3_cachedata_MPORT_data : _GEN_6834; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6836 = _GEN_8528 & 4'h4 == EntId[3:0] ? dataArray_42_4_cachedata_MPORT_data : _GEN_6835; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6837 = _GEN_8528 & 4'h5 == EntId[3:0] ? dataArray_42_5_cachedata_MPORT_data : _GEN_6836; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6838 = _GEN_8528 & 4'h6 == EntId[3:0] ? dataArray_42_6_cachedata_MPORT_data : _GEN_6837; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6839 = _GEN_8528 & 4'h7 == EntId[3:0] ? dataArray_42_7_cachedata_MPORT_data : _GEN_6838; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6840 = _GEN_8528 & 4'h8 == EntId[3:0] ? dataArray_42_8_cachedata_MPORT_data : _GEN_6839; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6841 = _GEN_8528 & 4'h9 == EntId[3:0] ? dataArray_42_9_cachedata_MPORT_data : _GEN_6840; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6842 = _GEN_8528 & 4'ha == EntId[3:0] ? dataArray_42_10_cachedata_MPORT_data : _GEN_6841; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6843 = _GEN_8528 & 4'hb == EntId[3:0] ? dataArray_42_11_cachedata_MPORT_data : _GEN_6842; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6844 = _GEN_8528 & 4'hc == EntId[3:0] ? dataArray_42_12_cachedata_MPORT_data : _GEN_6843; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6845 = _GEN_8528 & 4'hd == EntId[3:0] ? dataArray_42_13_cachedata_MPORT_data : _GEN_6844; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6846 = _GEN_8528 & 4'he == EntId[3:0] ? dataArray_42_14_cachedata_MPORT_data : _GEN_6845; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6847 = _GEN_8528 & 4'hf == EntId[3:0] ? dataArray_42_15_cachedata_MPORT_data : _GEN_6846; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6848 = _GEN_8560 & 4'h0 == EntId[3:0] ? dataArray_43_0_cachedata_MPORT_data : _GEN_6847; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6849 = _GEN_8560 & 4'h1 == EntId[3:0] ? dataArray_43_1_cachedata_MPORT_data : _GEN_6848; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6850 = _GEN_8560 & 4'h2 == EntId[3:0] ? dataArray_43_2_cachedata_MPORT_data : _GEN_6849; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6851 = _GEN_8560 & 4'h3 == EntId[3:0] ? dataArray_43_3_cachedata_MPORT_data : _GEN_6850; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6852 = _GEN_8560 & 4'h4 == EntId[3:0] ? dataArray_43_4_cachedata_MPORT_data : _GEN_6851; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6853 = _GEN_8560 & 4'h5 == EntId[3:0] ? dataArray_43_5_cachedata_MPORT_data : _GEN_6852; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6854 = _GEN_8560 & 4'h6 == EntId[3:0] ? dataArray_43_6_cachedata_MPORT_data : _GEN_6853; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6855 = _GEN_8560 & 4'h7 == EntId[3:0] ? dataArray_43_7_cachedata_MPORT_data : _GEN_6854; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6856 = _GEN_8560 & 4'h8 == EntId[3:0] ? dataArray_43_8_cachedata_MPORT_data : _GEN_6855; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6857 = _GEN_8560 & 4'h9 == EntId[3:0] ? dataArray_43_9_cachedata_MPORT_data : _GEN_6856; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6858 = _GEN_8560 & 4'ha == EntId[3:0] ? dataArray_43_10_cachedata_MPORT_data : _GEN_6857; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6859 = _GEN_8560 & 4'hb == EntId[3:0] ? dataArray_43_11_cachedata_MPORT_data : _GEN_6858; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6860 = _GEN_8560 & 4'hc == EntId[3:0] ? dataArray_43_12_cachedata_MPORT_data : _GEN_6859; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6861 = _GEN_8560 & 4'hd == EntId[3:0] ? dataArray_43_13_cachedata_MPORT_data : _GEN_6860; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6862 = _GEN_8560 & 4'he == EntId[3:0] ? dataArray_43_14_cachedata_MPORT_data : _GEN_6861; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6863 = _GEN_8560 & 4'hf == EntId[3:0] ? dataArray_43_15_cachedata_MPORT_data : _GEN_6862; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6864 = _GEN_8592 & 4'h0 == EntId[3:0] ? dataArray_44_0_cachedata_MPORT_data : _GEN_6863; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6865 = _GEN_8592 & 4'h1 == EntId[3:0] ? dataArray_44_1_cachedata_MPORT_data : _GEN_6864; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6866 = _GEN_8592 & 4'h2 == EntId[3:0] ? dataArray_44_2_cachedata_MPORT_data : _GEN_6865; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6867 = _GEN_8592 & 4'h3 == EntId[3:0] ? dataArray_44_3_cachedata_MPORT_data : _GEN_6866; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6868 = _GEN_8592 & 4'h4 == EntId[3:0] ? dataArray_44_4_cachedata_MPORT_data : _GEN_6867; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6869 = _GEN_8592 & 4'h5 == EntId[3:0] ? dataArray_44_5_cachedata_MPORT_data : _GEN_6868; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6870 = _GEN_8592 & 4'h6 == EntId[3:0] ? dataArray_44_6_cachedata_MPORT_data : _GEN_6869; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6871 = _GEN_8592 & 4'h7 == EntId[3:0] ? dataArray_44_7_cachedata_MPORT_data : _GEN_6870; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6872 = _GEN_8592 & 4'h8 == EntId[3:0] ? dataArray_44_8_cachedata_MPORT_data : _GEN_6871; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6873 = _GEN_8592 & 4'h9 == EntId[3:0] ? dataArray_44_9_cachedata_MPORT_data : _GEN_6872; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6874 = _GEN_8592 & 4'ha == EntId[3:0] ? dataArray_44_10_cachedata_MPORT_data : _GEN_6873; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6875 = _GEN_8592 & 4'hb == EntId[3:0] ? dataArray_44_11_cachedata_MPORT_data : _GEN_6874; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6876 = _GEN_8592 & 4'hc == EntId[3:0] ? dataArray_44_12_cachedata_MPORT_data : _GEN_6875; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6877 = _GEN_8592 & 4'hd == EntId[3:0] ? dataArray_44_13_cachedata_MPORT_data : _GEN_6876; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6878 = _GEN_8592 & 4'he == EntId[3:0] ? dataArray_44_14_cachedata_MPORT_data : _GEN_6877; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6879 = _GEN_8592 & 4'hf == EntId[3:0] ? dataArray_44_15_cachedata_MPORT_data : _GEN_6878; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6880 = _GEN_8624 & 4'h0 == EntId[3:0] ? dataArray_45_0_cachedata_MPORT_data : _GEN_6879; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6881 = _GEN_8624 & 4'h1 == EntId[3:0] ? dataArray_45_1_cachedata_MPORT_data : _GEN_6880; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6882 = _GEN_8624 & 4'h2 == EntId[3:0] ? dataArray_45_2_cachedata_MPORT_data : _GEN_6881; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6883 = _GEN_8624 & 4'h3 == EntId[3:0] ? dataArray_45_3_cachedata_MPORT_data : _GEN_6882; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6884 = _GEN_8624 & 4'h4 == EntId[3:0] ? dataArray_45_4_cachedata_MPORT_data : _GEN_6883; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6885 = _GEN_8624 & 4'h5 == EntId[3:0] ? dataArray_45_5_cachedata_MPORT_data : _GEN_6884; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6886 = _GEN_8624 & 4'h6 == EntId[3:0] ? dataArray_45_6_cachedata_MPORT_data : _GEN_6885; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6887 = _GEN_8624 & 4'h7 == EntId[3:0] ? dataArray_45_7_cachedata_MPORT_data : _GEN_6886; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6888 = _GEN_8624 & 4'h8 == EntId[3:0] ? dataArray_45_8_cachedata_MPORT_data : _GEN_6887; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6889 = _GEN_8624 & 4'h9 == EntId[3:0] ? dataArray_45_9_cachedata_MPORT_data : _GEN_6888; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6890 = _GEN_8624 & 4'ha == EntId[3:0] ? dataArray_45_10_cachedata_MPORT_data : _GEN_6889; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6891 = _GEN_8624 & 4'hb == EntId[3:0] ? dataArray_45_11_cachedata_MPORT_data : _GEN_6890; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6892 = _GEN_8624 & 4'hc == EntId[3:0] ? dataArray_45_12_cachedata_MPORT_data : _GEN_6891; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6893 = _GEN_8624 & 4'hd == EntId[3:0] ? dataArray_45_13_cachedata_MPORT_data : _GEN_6892; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6894 = _GEN_8624 & 4'he == EntId[3:0] ? dataArray_45_14_cachedata_MPORT_data : _GEN_6893; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6895 = _GEN_8624 & 4'hf == EntId[3:0] ? dataArray_45_15_cachedata_MPORT_data : _GEN_6894; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6896 = _GEN_8656 & 4'h0 == EntId[3:0] ? dataArray_46_0_cachedata_MPORT_data : _GEN_6895; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6897 = _GEN_8656 & 4'h1 == EntId[3:0] ? dataArray_46_1_cachedata_MPORT_data : _GEN_6896; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6898 = _GEN_8656 & 4'h2 == EntId[3:0] ? dataArray_46_2_cachedata_MPORT_data : _GEN_6897; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6899 = _GEN_8656 & 4'h3 == EntId[3:0] ? dataArray_46_3_cachedata_MPORT_data : _GEN_6898; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6900 = _GEN_8656 & 4'h4 == EntId[3:0] ? dataArray_46_4_cachedata_MPORT_data : _GEN_6899; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6901 = _GEN_8656 & 4'h5 == EntId[3:0] ? dataArray_46_5_cachedata_MPORT_data : _GEN_6900; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6902 = _GEN_8656 & 4'h6 == EntId[3:0] ? dataArray_46_6_cachedata_MPORT_data : _GEN_6901; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6903 = _GEN_8656 & 4'h7 == EntId[3:0] ? dataArray_46_7_cachedata_MPORT_data : _GEN_6902; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6904 = _GEN_8656 & 4'h8 == EntId[3:0] ? dataArray_46_8_cachedata_MPORT_data : _GEN_6903; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6905 = _GEN_8656 & 4'h9 == EntId[3:0] ? dataArray_46_9_cachedata_MPORT_data : _GEN_6904; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6906 = _GEN_8656 & 4'ha == EntId[3:0] ? dataArray_46_10_cachedata_MPORT_data : _GEN_6905; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6907 = _GEN_8656 & 4'hb == EntId[3:0] ? dataArray_46_11_cachedata_MPORT_data : _GEN_6906; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6908 = _GEN_8656 & 4'hc == EntId[3:0] ? dataArray_46_12_cachedata_MPORT_data : _GEN_6907; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6909 = _GEN_8656 & 4'hd == EntId[3:0] ? dataArray_46_13_cachedata_MPORT_data : _GEN_6908; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6910 = _GEN_8656 & 4'he == EntId[3:0] ? dataArray_46_14_cachedata_MPORT_data : _GEN_6909; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6911 = _GEN_8656 & 4'hf == EntId[3:0] ? dataArray_46_15_cachedata_MPORT_data : _GEN_6910; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6912 = _GEN_8688 & 4'h0 == EntId[3:0] ? dataArray_47_0_cachedata_MPORT_data : _GEN_6911; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6913 = _GEN_8688 & 4'h1 == EntId[3:0] ? dataArray_47_1_cachedata_MPORT_data : _GEN_6912; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6914 = _GEN_8688 & 4'h2 == EntId[3:0] ? dataArray_47_2_cachedata_MPORT_data : _GEN_6913; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6915 = _GEN_8688 & 4'h3 == EntId[3:0] ? dataArray_47_3_cachedata_MPORT_data : _GEN_6914; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6916 = _GEN_8688 & 4'h4 == EntId[3:0] ? dataArray_47_4_cachedata_MPORT_data : _GEN_6915; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6917 = _GEN_8688 & 4'h5 == EntId[3:0] ? dataArray_47_5_cachedata_MPORT_data : _GEN_6916; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6918 = _GEN_8688 & 4'h6 == EntId[3:0] ? dataArray_47_6_cachedata_MPORT_data : _GEN_6917; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6919 = _GEN_8688 & 4'h7 == EntId[3:0] ? dataArray_47_7_cachedata_MPORT_data : _GEN_6918; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6920 = _GEN_8688 & 4'h8 == EntId[3:0] ? dataArray_47_8_cachedata_MPORT_data : _GEN_6919; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6921 = _GEN_8688 & 4'h9 == EntId[3:0] ? dataArray_47_9_cachedata_MPORT_data : _GEN_6920; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6922 = _GEN_8688 & 4'ha == EntId[3:0] ? dataArray_47_10_cachedata_MPORT_data : _GEN_6921; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6923 = _GEN_8688 & 4'hb == EntId[3:0] ? dataArray_47_11_cachedata_MPORT_data : _GEN_6922; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6924 = _GEN_8688 & 4'hc == EntId[3:0] ? dataArray_47_12_cachedata_MPORT_data : _GEN_6923; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6925 = _GEN_8688 & 4'hd == EntId[3:0] ? dataArray_47_13_cachedata_MPORT_data : _GEN_6924; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6926 = _GEN_8688 & 4'he == EntId[3:0] ? dataArray_47_14_cachedata_MPORT_data : _GEN_6925; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6927 = _GEN_8688 & 4'hf == EntId[3:0] ? dataArray_47_15_cachedata_MPORT_data : _GEN_6926; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6928 = _GEN_8720 & 4'h0 == EntId[3:0] ? dataArray_48_0_cachedata_MPORT_data : _GEN_6927; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6929 = _GEN_8720 & 4'h1 == EntId[3:0] ? dataArray_48_1_cachedata_MPORT_data : _GEN_6928; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6930 = _GEN_8720 & 4'h2 == EntId[3:0] ? dataArray_48_2_cachedata_MPORT_data : _GEN_6929; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6931 = _GEN_8720 & 4'h3 == EntId[3:0] ? dataArray_48_3_cachedata_MPORT_data : _GEN_6930; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6932 = _GEN_8720 & 4'h4 == EntId[3:0] ? dataArray_48_4_cachedata_MPORT_data : _GEN_6931; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6933 = _GEN_8720 & 4'h5 == EntId[3:0] ? dataArray_48_5_cachedata_MPORT_data : _GEN_6932; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6934 = _GEN_8720 & 4'h6 == EntId[3:0] ? dataArray_48_6_cachedata_MPORT_data : _GEN_6933; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6935 = _GEN_8720 & 4'h7 == EntId[3:0] ? dataArray_48_7_cachedata_MPORT_data : _GEN_6934; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6936 = _GEN_8720 & 4'h8 == EntId[3:0] ? dataArray_48_8_cachedata_MPORT_data : _GEN_6935; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6937 = _GEN_8720 & 4'h9 == EntId[3:0] ? dataArray_48_9_cachedata_MPORT_data : _GEN_6936; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6938 = _GEN_8720 & 4'ha == EntId[3:0] ? dataArray_48_10_cachedata_MPORT_data : _GEN_6937; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6939 = _GEN_8720 & 4'hb == EntId[3:0] ? dataArray_48_11_cachedata_MPORT_data : _GEN_6938; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6940 = _GEN_8720 & 4'hc == EntId[3:0] ? dataArray_48_12_cachedata_MPORT_data : _GEN_6939; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6941 = _GEN_8720 & 4'hd == EntId[3:0] ? dataArray_48_13_cachedata_MPORT_data : _GEN_6940; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6942 = _GEN_8720 & 4'he == EntId[3:0] ? dataArray_48_14_cachedata_MPORT_data : _GEN_6941; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6943 = _GEN_8720 & 4'hf == EntId[3:0] ? dataArray_48_15_cachedata_MPORT_data : _GEN_6942; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6944 = _GEN_8752 & 4'h0 == EntId[3:0] ? dataArray_49_0_cachedata_MPORT_data : _GEN_6943; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6945 = _GEN_8752 & 4'h1 == EntId[3:0] ? dataArray_49_1_cachedata_MPORT_data : _GEN_6944; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6946 = _GEN_8752 & 4'h2 == EntId[3:0] ? dataArray_49_2_cachedata_MPORT_data : _GEN_6945; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6947 = _GEN_8752 & 4'h3 == EntId[3:0] ? dataArray_49_3_cachedata_MPORT_data : _GEN_6946; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6948 = _GEN_8752 & 4'h4 == EntId[3:0] ? dataArray_49_4_cachedata_MPORT_data : _GEN_6947; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6949 = _GEN_8752 & 4'h5 == EntId[3:0] ? dataArray_49_5_cachedata_MPORT_data : _GEN_6948; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6950 = _GEN_8752 & 4'h6 == EntId[3:0] ? dataArray_49_6_cachedata_MPORT_data : _GEN_6949; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6951 = _GEN_8752 & 4'h7 == EntId[3:0] ? dataArray_49_7_cachedata_MPORT_data : _GEN_6950; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6952 = _GEN_8752 & 4'h8 == EntId[3:0] ? dataArray_49_8_cachedata_MPORT_data : _GEN_6951; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6953 = _GEN_8752 & 4'h9 == EntId[3:0] ? dataArray_49_9_cachedata_MPORT_data : _GEN_6952; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6954 = _GEN_8752 & 4'ha == EntId[3:0] ? dataArray_49_10_cachedata_MPORT_data : _GEN_6953; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6955 = _GEN_8752 & 4'hb == EntId[3:0] ? dataArray_49_11_cachedata_MPORT_data : _GEN_6954; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6956 = _GEN_8752 & 4'hc == EntId[3:0] ? dataArray_49_12_cachedata_MPORT_data : _GEN_6955; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6957 = _GEN_8752 & 4'hd == EntId[3:0] ? dataArray_49_13_cachedata_MPORT_data : _GEN_6956; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6958 = _GEN_8752 & 4'he == EntId[3:0] ? dataArray_49_14_cachedata_MPORT_data : _GEN_6957; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6959 = _GEN_8752 & 4'hf == EntId[3:0] ? dataArray_49_15_cachedata_MPORT_data : _GEN_6958; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6960 = _GEN_8784 & 4'h0 == EntId[3:0] ? dataArray_50_0_cachedata_MPORT_data : _GEN_6959; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6961 = _GEN_8784 & 4'h1 == EntId[3:0] ? dataArray_50_1_cachedata_MPORT_data : _GEN_6960; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6962 = _GEN_8784 & 4'h2 == EntId[3:0] ? dataArray_50_2_cachedata_MPORT_data : _GEN_6961; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6963 = _GEN_8784 & 4'h3 == EntId[3:0] ? dataArray_50_3_cachedata_MPORT_data : _GEN_6962; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6964 = _GEN_8784 & 4'h4 == EntId[3:0] ? dataArray_50_4_cachedata_MPORT_data : _GEN_6963; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6965 = _GEN_8784 & 4'h5 == EntId[3:0] ? dataArray_50_5_cachedata_MPORT_data : _GEN_6964; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6966 = _GEN_8784 & 4'h6 == EntId[3:0] ? dataArray_50_6_cachedata_MPORT_data : _GEN_6965; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6967 = _GEN_8784 & 4'h7 == EntId[3:0] ? dataArray_50_7_cachedata_MPORT_data : _GEN_6966; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6968 = _GEN_8784 & 4'h8 == EntId[3:0] ? dataArray_50_8_cachedata_MPORT_data : _GEN_6967; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6969 = _GEN_8784 & 4'h9 == EntId[3:0] ? dataArray_50_9_cachedata_MPORT_data : _GEN_6968; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6970 = _GEN_8784 & 4'ha == EntId[3:0] ? dataArray_50_10_cachedata_MPORT_data : _GEN_6969; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6971 = _GEN_8784 & 4'hb == EntId[3:0] ? dataArray_50_11_cachedata_MPORT_data : _GEN_6970; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6972 = _GEN_8784 & 4'hc == EntId[3:0] ? dataArray_50_12_cachedata_MPORT_data : _GEN_6971; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6973 = _GEN_8784 & 4'hd == EntId[3:0] ? dataArray_50_13_cachedata_MPORT_data : _GEN_6972; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6974 = _GEN_8784 & 4'he == EntId[3:0] ? dataArray_50_14_cachedata_MPORT_data : _GEN_6973; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6975 = _GEN_8784 & 4'hf == EntId[3:0] ? dataArray_50_15_cachedata_MPORT_data : _GEN_6974; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6976 = _GEN_8816 & 4'h0 == EntId[3:0] ? dataArray_51_0_cachedata_MPORT_data : _GEN_6975; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6977 = _GEN_8816 & 4'h1 == EntId[3:0] ? dataArray_51_1_cachedata_MPORT_data : _GEN_6976; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6978 = _GEN_8816 & 4'h2 == EntId[3:0] ? dataArray_51_2_cachedata_MPORT_data : _GEN_6977; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6979 = _GEN_8816 & 4'h3 == EntId[3:0] ? dataArray_51_3_cachedata_MPORT_data : _GEN_6978; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6980 = _GEN_8816 & 4'h4 == EntId[3:0] ? dataArray_51_4_cachedata_MPORT_data : _GEN_6979; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6981 = _GEN_8816 & 4'h5 == EntId[3:0] ? dataArray_51_5_cachedata_MPORT_data : _GEN_6980; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6982 = _GEN_8816 & 4'h6 == EntId[3:0] ? dataArray_51_6_cachedata_MPORT_data : _GEN_6981; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6983 = _GEN_8816 & 4'h7 == EntId[3:0] ? dataArray_51_7_cachedata_MPORT_data : _GEN_6982; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6984 = _GEN_8816 & 4'h8 == EntId[3:0] ? dataArray_51_8_cachedata_MPORT_data : _GEN_6983; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6985 = _GEN_8816 & 4'h9 == EntId[3:0] ? dataArray_51_9_cachedata_MPORT_data : _GEN_6984; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6986 = _GEN_8816 & 4'ha == EntId[3:0] ? dataArray_51_10_cachedata_MPORT_data : _GEN_6985; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6987 = _GEN_8816 & 4'hb == EntId[3:0] ? dataArray_51_11_cachedata_MPORT_data : _GEN_6986; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6988 = _GEN_8816 & 4'hc == EntId[3:0] ? dataArray_51_12_cachedata_MPORT_data : _GEN_6987; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6989 = _GEN_8816 & 4'hd == EntId[3:0] ? dataArray_51_13_cachedata_MPORT_data : _GEN_6988; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6990 = _GEN_8816 & 4'he == EntId[3:0] ? dataArray_51_14_cachedata_MPORT_data : _GEN_6989; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6991 = _GEN_8816 & 4'hf == EntId[3:0] ? dataArray_51_15_cachedata_MPORT_data : _GEN_6990; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6992 = _GEN_8848 & 4'h0 == EntId[3:0] ? dataArray_52_0_cachedata_MPORT_data : _GEN_6991; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6993 = _GEN_8848 & 4'h1 == EntId[3:0] ? dataArray_52_1_cachedata_MPORT_data : _GEN_6992; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6994 = _GEN_8848 & 4'h2 == EntId[3:0] ? dataArray_52_2_cachedata_MPORT_data : _GEN_6993; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6995 = _GEN_8848 & 4'h3 == EntId[3:0] ? dataArray_52_3_cachedata_MPORT_data : _GEN_6994; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6996 = _GEN_8848 & 4'h4 == EntId[3:0] ? dataArray_52_4_cachedata_MPORT_data : _GEN_6995; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6997 = _GEN_8848 & 4'h5 == EntId[3:0] ? dataArray_52_5_cachedata_MPORT_data : _GEN_6996; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6998 = _GEN_8848 & 4'h6 == EntId[3:0] ? dataArray_52_6_cachedata_MPORT_data : _GEN_6997; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_6999 = _GEN_8848 & 4'h7 == EntId[3:0] ? dataArray_52_7_cachedata_MPORT_data : _GEN_6998; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7000 = _GEN_8848 & 4'h8 == EntId[3:0] ? dataArray_52_8_cachedata_MPORT_data : _GEN_6999; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7001 = _GEN_8848 & 4'h9 == EntId[3:0] ? dataArray_52_9_cachedata_MPORT_data : _GEN_7000; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7002 = _GEN_8848 & 4'ha == EntId[3:0] ? dataArray_52_10_cachedata_MPORT_data : _GEN_7001; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7003 = _GEN_8848 & 4'hb == EntId[3:0] ? dataArray_52_11_cachedata_MPORT_data : _GEN_7002; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7004 = _GEN_8848 & 4'hc == EntId[3:0] ? dataArray_52_12_cachedata_MPORT_data : _GEN_7003; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7005 = _GEN_8848 & 4'hd == EntId[3:0] ? dataArray_52_13_cachedata_MPORT_data : _GEN_7004; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7006 = _GEN_8848 & 4'he == EntId[3:0] ? dataArray_52_14_cachedata_MPORT_data : _GEN_7005; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7007 = _GEN_8848 & 4'hf == EntId[3:0] ? dataArray_52_15_cachedata_MPORT_data : _GEN_7006; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7008 = _GEN_8880 & 4'h0 == EntId[3:0] ? dataArray_53_0_cachedata_MPORT_data : _GEN_7007; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7009 = _GEN_8880 & 4'h1 == EntId[3:0] ? dataArray_53_1_cachedata_MPORT_data : _GEN_7008; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7010 = _GEN_8880 & 4'h2 == EntId[3:0] ? dataArray_53_2_cachedata_MPORT_data : _GEN_7009; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7011 = _GEN_8880 & 4'h3 == EntId[3:0] ? dataArray_53_3_cachedata_MPORT_data : _GEN_7010; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7012 = _GEN_8880 & 4'h4 == EntId[3:0] ? dataArray_53_4_cachedata_MPORT_data : _GEN_7011; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7013 = _GEN_8880 & 4'h5 == EntId[3:0] ? dataArray_53_5_cachedata_MPORT_data : _GEN_7012; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7014 = _GEN_8880 & 4'h6 == EntId[3:0] ? dataArray_53_6_cachedata_MPORT_data : _GEN_7013; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7015 = _GEN_8880 & 4'h7 == EntId[3:0] ? dataArray_53_7_cachedata_MPORT_data : _GEN_7014; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7016 = _GEN_8880 & 4'h8 == EntId[3:0] ? dataArray_53_8_cachedata_MPORT_data : _GEN_7015; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7017 = _GEN_8880 & 4'h9 == EntId[3:0] ? dataArray_53_9_cachedata_MPORT_data : _GEN_7016; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7018 = _GEN_8880 & 4'ha == EntId[3:0] ? dataArray_53_10_cachedata_MPORT_data : _GEN_7017; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7019 = _GEN_8880 & 4'hb == EntId[3:0] ? dataArray_53_11_cachedata_MPORT_data : _GEN_7018; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7020 = _GEN_8880 & 4'hc == EntId[3:0] ? dataArray_53_12_cachedata_MPORT_data : _GEN_7019; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7021 = _GEN_8880 & 4'hd == EntId[3:0] ? dataArray_53_13_cachedata_MPORT_data : _GEN_7020; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7022 = _GEN_8880 & 4'he == EntId[3:0] ? dataArray_53_14_cachedata_MPORT_data : _GEN_7021; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7023 = _GEN_8880 & 4'hf == EntId[3:0] ? dataArray_53_15_cachedata_MPORT_data : _GEN_7022; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7024 = _GEN_8912 & 4'h0 == EntId[3:0] ? dataArray_54_0_cachedata_MPORT_data : _GEN_7023; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7025 = _GEN_8912 & 4'h1 == EntId[3:0] ? dataArray_54_1_cachedata_MPORT_data : _GEN_7024; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7026 = _GEN_8912 & 4'h2 == EntId[3:0] ? dataArray_54_2_cachedata_MPORT_data : _GEN_7025; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7027 = _GEN_8912 & 4'h3 == EntId[3:0] ? dataArray_54_3_cachedata_MPORT_data : _GEN_7026; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7028 = _GEN_8912 & 4'h4 == EntId[3:0] ? dataArray_54_4_cachedata_MPORT_data : _GEN_7027; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7029 = _GEN_8912 & 4'h5 == EntId[3:0] ? dataArray_54_5_cachedata_MPORT_data : _GEN_7028; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7030 = _GEN_8912 & 4'h6 == EntId[3:0] ? dataArray_54_6_cachedata_MPORT_data : _GEN_7029; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7031 = _GEN_8912 & 4'h7 == EntId[3:0] ? dataArray_54_7_cachedata_MPORT_data : _GEN_7030; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7032 = _GEN_8912 & 4'h8 == EntId[3:0] ? dataArray_54_8_cachedata_MPORT_data : _GEN_7031; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7033 = _GEN_8912 & 4'h9 == EntId[3:0] ? dataArray_54_9_cachedata_MPORT_data : _GEN_7032; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7034 = _GEN_8912 & 4'ha == EntId[3:0] ? dataArray_54_10_cachedata_MPORT_data : _GEN_7033; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7035 = _GEN_8912 & 4'hb == EntId[3:0] ? dataArray_54_11_cachedata_MPORT_data : _GEN_7034; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7036 = _GEN_8912 & 4'hc == EntId[3:0] ? dataArray_54_12_cachedata_MPORT_data : _GEN_7035; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7037 = _GEN_8912 & 4'hd == EntId[3:0] ? dataArray_54_13_cachedata_MPORT_data : _GEN_7036; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7038 = _GEN_8912 & 4'he == EntId[3:0] ? dataArray_54_14_cachedata_MPORT_data : _GEN_7037; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7039 = _GEN_8912 & 4'hf == EntId[3:0] ? dataArray_54_15_cachedata_MPORT_data : _GEN_7038; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7040 = _GEN_8944 & 4'h0 == EntId[3:0] ? dataArray_55_0_cachedata_MPORT_data : _GEN_7039; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7041 = _GEN_8944 & 4'h1 == EntId[3:0] ? dataArray_55_1_cachedata_MPORT_data : _GEN_7040; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7042 = _GEN_8944 & 4'h2 == EntId[3:0] ? dataArray_55_2_cachedata_MPORT_data : _GEN_7041; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7043 = _GEN_8944 & 4'h3 == EntId[3:0] ? dataArray_55_3_cachedata_MPORT_data : _GEN_7042; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7044 = _GEN_8944 & 4'h4 == EntId[3:0] ? dataArray_55_4_cachedata_MPORT_data : _GEN_7043; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7045 = _GEN_8944 & 4'h5 == EntId[3:0] ? dataArray_55_5_cachedata_MPORT_data : _GEN_7044; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7046 = _GEN_8944 & 4'h6 == EntId[3:0] ? dataArray_55_6_cachedata_MPORT_data : _GEN_7045; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7047 = _GEN_8944 & 4'h7 == EntId[3:0] ? dataArray_55_7_cachedata_MPORT_data : _GEN_7046; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7048 = _GEN_8944 & 4'h8 == EntId[3:0] ? dataArray_55_8_cachedata_MPORT_data : _GEN_7047; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7049 = _GEN_8944 & 4'h9 == EntId[3:0] ? dataArray_55_9_cachedata_MPORT_data : _GEN_7048; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7050 = _GEN_8944 & 4'ha == EntId[3:0] ? dataArray_55_10_cachedata_MPORT_data : _GEN_7049; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7051 = _GEN_8944 & 4'hb == EntId[3:0] ? dataArray_55_11_cachedata_MPORT_data : _GEN_7050; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7052 = _GEN_8944 & 4'hc == EntId[3:0] ? dataArray_55_12_cachedata_MPORT_data : _GEN_7051; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7053 = _GEN_8944 & 4'hd == EntId[3:0] ? dataArray_55_13_cachedata_MPORT_data : _GEN_7052; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7054 = _GEN_8944 & 4'he == EntId[3:0] ? dataArray_55_14_cachedata_MPORT_data : _GEN_7053; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7055 = _GEN_8944 & 4'hf == EntId[3:0] ? dataArray_55_15_cachedata_MPORT_data : _GEN_7054; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7056 = _GEN_8976 & 4'h0 == EntId[3:0] ? dataArray_56_0_cachedata_MPORT_data : _GEN_7055; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7057 = _GEN_8976 & 4'h1 == EntId[3:0] ? dataArray_56_1_cachedata_MPORT_data : _GEN_7056; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7058 = _GEN_8976 & 4'h2 == EntId[3:0] ? dataArray_56_2_cachedata_MPORT_data : _GEN_7057; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7059 = _GEN_8976 & 4'h3 == EntId[3:0] ? dataArray_56_3_cachedata_MPORT_data : _GEN_7058; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7060 = _GEN_8976 & 4'h4 == EntId[3:0] ? dataArray_56_4_cachedata_MPORT_data : _GEN_7059; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7061 = _GEN_8976 & 4'h5 == EntId[3:0] ? dataArray_56_5_cachedata_MPORT_data : _GEN_7060; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7062 = _GEN_8976 & 4'h6 == EntId[3:0] ? dataArray_56_6_cachedata_MPORT_data : _GEN_7061; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7063 = _GEN_8976 & 4'h7 == EntId[3:0] ? dataArray_56_7_cachedata_MPORT_data : _GEN_7062; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7064 = _GEN_8976 & 4'h8 == EntId[3:0] ? dataArray_56_8_cachedata_MPORT_data : _GEN_7063; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7065 = _GEN_8976 & 4'h9 == EntId[3:0] ? dataArray_56_9_cachedata_MPORT_data : _GEN_7064; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7066 = _GEN_8976 & 4'ha == EntId[3:0] ? dataArray_56_10_cachedata_MPORT_data : _GEN_7065; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7067 = _GEN_8976 & 4'hb == EntId[3:0] ? dataArray_56_11_cachedata_MPORT_data : _GEN_7066; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7068 = _GEN_8976 & 4'hc == EntId[3:0] ? dataArray_56_12_cachedata_MPORT_data : _GEN_7067; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7069 = _GEN_8976 & 4'hd == EntId[3:0] ? dataArray_56_13_cachedata_MPORT_data : _GEN_7068; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7070 = _GEN_8976 & 4'he == EntId[3:0] ? dataArray_56_14_cachedata_MPORT_data : _GEN_7069; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7071 = _GEN_8976 & 4'hf == EntId[3:0] ? dataArray_56_15_cachedata_MPORT_data : _GEN_7070; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7072 = _GEN_9008 & 4'h0 == EntId[3:0] ? dataArray_57_0_cachedata_MPORT_data : _GEN_7071; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7073 = _GEN_9008 & 4'h1 == EntId[3:0] ? dataArray_57_1_cachedata_MPORT_data : _GEN_7072; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7074 = _GEN_9008 & 4'h2 == EntId[3:0] ? dataArray_57_2_cachedata_MPORT_data : _GEN_7073; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7075 = _GEN_9008 & 4'h3 == EntId[3:0] ? dataArray_57_3_cachedata_MPORT_data : _GEN_7074; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7076 = _GEN_9008 & 4'h4 == EntId[3:0] ? dataArray_57_4_cachedata_MPORT_data : _GEN_7075; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7077 = _GEN_9008 & 4'h5 == EntId[3:0] ? dataArray_57_5_cachedata_MPORT_data : _GEN_7076; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7078 = _GEN_9008 & 4'h6 == EntId[3:0] ? dataArray_57_6_cachedata_MPORT_data : _GEN_7077; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7079 = _GEN_9008 & 4'h7 == EntId[3:0] ? dataArray_57_7_cachedata_MPORT_data : _GEN_7078; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7080 = _GEN_9008 & 4'h8 == EntId[3:0] ? dataArray_57_8_cachedata_MPORT_data : _GEN_7079; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7081 = _GEN_9008 & 4'h9 == EntId[3:0] ? dataArray_57_9_cachedata_MPORT_data : _GEN_7080; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7082 = _GEN_9008 & 4'ha == EntId[3:0] ? dataArray_57_10_cachedata_MPORT_data : _GEN_7081; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7083 = _GEN_9008 & 4'hb == EntId[3:0] ? dataArray_57_11_cachedata_MPORT_data : _GEN_7082; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7084 = _GEN_9008 & 4'hc == EntId[3:0] ? dataArray_57_12_cachedata_MPORT_data : _GEN_7083; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7085 = _GEN_9008 & 4'hd == EntId[3:0] ? dataArray_57_13_cachedata_MPORT_data : _GEN_7084; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7086 = _GEN_9008 & 4'he == EntId[3:0] ? dataArray_57_14_cachedata_MPORT_data : _GEN_7085; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7087 = _GEN_9008 & 4'hf == EntId[3:0] ? dataArray_57_15_cachedata_MPORT_data : _GEN_7086; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7088 = _GEN_9040 & 4'h0 == EntId[3:0] ? dataArray_58_0_cachedata_MPORT_data : _GEN_7087; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7089 = _GEN_9040 & 4'h1 == EntId[3:0] ? dataArray_58_1_cachedata_MPORT_data : _GEN_7088; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7090 = _GEN_9040 & 4'h2 == EntId[3:0] ? dataArray_58_2_cachedata_MPORT_data : _GEN_7089; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7091 = _GEN_9040 & 4'h3 == EntId[3:0] ? dataArray_58_3_cachedata_MPORT_data : _GEN_7090; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7092 = _GEN_9040 & 4'h4 == EntId[3:0] ? dataArray_58_4_cachedata_MPORT_data : _GEN_7091; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7093 = _GEN_9040 & 4'h5 == EntId[3:0] ? dataArray_58_5_cachedata_MPORT_data : _GEN_7092; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7094 = _GEN_9040 & 4'h6 == EntId[3:0] ? dataArray_58_6_cachedata_MPORT_data : _GEN_7093; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7095 = _GEN_9040 & 4'h7 == EntId[3:0] ? dataArray_58_7_cachedata_MPORT_data : _GEN_7094; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7096 = _GEN_9040 & 4'h8 == EntId[3:0] ? dataArray_58_8_cachedata_MPORT_data : _GEN_7095; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7097 = _GEN_9040 & 4'h9 == EntId[3:0] ? dataArray_58_9_cachedata_MPORT_data : _GEN_7096; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7098 = _GEN_9040 & 4'ha == EntId[3:0] ? dataArray_58_10_cachedata_MPORT_data : _GEN_7097; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7099 = _GEN_9040 & 4'hb == EntId[3:0] ? dataArray_58_11_cachedata_MPORT_data : _GEN_7098; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7100 = _GEN_9040 & 4'hc == EntId[3:0] ? dataArray_58_12_cachedata_MPORT_data : _GEN_7099; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7101 = _GEN_9040 & 4'hd == EntId[3:0] ? dataArray_58_13_cachedata_MPORT_data : _GEN_7100; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7102 = _GEN_9040 & 4'he == EntId[3:0] ? dataArray_58_14_cachedata_MPORT_data : _GEN_7101; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7103 = _GEN_9040 & 4'hf == EntId[3:0] ? dataArray_58_15_cachedata_MPORT_data : _GEN_7102; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7104 = _GEN_9072 & 4'h0 == EntId[3:0] ? dataArray_59_0_cachedata_MPORT_data : _GEN_7103; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7105 = _GEN_9072 & 4'h1 == EntId[3:0] ? dataArray_59_1_cachedata_MPORT_data : _GEN_7104; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7106 = _GEN_9072 & 4'h2 == EntId[3:0] ? dataArray_59_2_cachedata_MPORT_data : _GEN_7105; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7107 = _GEN_9072 & 4'h3 == EntId[3:0] ? dataArray_59_3_cachedata_MPORT_data : _GEN_7106; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7108 = _GEN_9072 & 4'h4 == EntId[3:0] ? dataArray_59_4_cachedata_MPORT_data : _GEN_7107; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7109 = _GEN_9072 & 4'h5 == EntId[3:0] ? dataArray_59_5_cachedata_MPORT_data : _GEN_7108; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7110 = _GEN_9072 & 4'h6 == EntId[3:0] ? dataArray_59_6_cachedata_MPORT_data : _GEN_7109; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7111 = _GEN_9072 & 4'h7 == EntId[3:0] ? dataArray_59_7_cachedata_MPORT_data : _GEN_7110; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7112 = _GEN_9072 & 4'h8 == EntId[3:0] ? dataArray_59_8_cachedata_MPORT_data : _GEN_7111; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7113 = _GEN_9072 & 4'h9 == EntId[3:0] ? dataArray_59_9_cachedata_MPORT_data : _GEN_7112; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7114 = _GEN_9072 & 4'ha == EntId[3:0] ? dataArray_59_10_cachedata_MPORT_data : _GEN_7113; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7115 = _GEN_9072 & 4'hb == EntId[3:0] ? dataArray_59_11_cachedata_MPORT_data : _GEN_7114; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7116 = _GEN_9072 & 4'hc == EntId[3:0] ? dataArray_59_12_cachedata_MPORT_data : _GEN_7115; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7117 = _GEN_9072 & 4'hd == EntId[3:0] ? dataArray_59_13_cachedata_MPORT_data : _GEN_7116; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7118 = _GEN_9072 & 4'he == EntId[3:0] ? dataArray_59_14_cachedata_MPORT_data : _GEN_7117; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7119 = _GEN_9072 & 4'hf == EntId[3:0] ? dataArray_59_15_cachedata_MPORT_data : _GEN_7118; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7120 = _GEN_9104 & 4'h0 == EntId[3:0] ? dataArray_60_0_cachedata_MPORT_data : _GEN_7119; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7121 = _GEN_9104 & 4'h1 == EntId[3:0] ? dataArray_60_1_cachedata_MPORT_data : _GEN_7120; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7122 = _GEN_9104 & 4'h2 == EntId[3:0] ? dataArray_60_2_cachedata_MPORT_data : _GEN_7121; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7123 = _GEN_9104 & 4'h3 == EntId[3:0] ? dataArray_60_3_cachedata_MPORT_data : _GEN_7122; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7124 = _GEN_9104 & 4'h4 == EntId[3:0] ? dataArray_60_4_cachedata_MPORT_data : _GEN_7123; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7125 = _GEN_9104 & 4'h5 == EntId[3:0] ? dataArray_60_5_cachedata_MPORT_data : _GEN_7124; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7126 = _GEN_9104 & 4'h6 == EntId[3:0] ? dataArray_60_6_cachedata_MPORT_data : _GEN_7125; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7127 = _GEN_9104 & 4'h7 == EntId[3:0] ? dataArray_60_7_cachedata_MPORT_data : _GEN_7126; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7128 = _GEN_9104 & 4'h8 == EntId[3:0] ? dataArray_60_8_cachedata_MPORT_data : _GEN_7127; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7129 = _GEN_9104 & 4'h9 == EntId[3:0] ? dataArray_60_9_cachedata_MPORT_data : _GEN_7128; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7130 = _GEN_9104 & 4'ha == EntId[3:0] ? dataArray_60_10_cachedata_MPORT_data : _GEN_7129; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7131 = _GEN_9104 & 4'hb == EntId[3:0] ? dataArray_60_11_cachedata_MPORT_data : _GEN_7130; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7132 = _GEN_9104 & 4'hc == EntId[3:0] ? dataArray_60_12_cachedata_MPORT_data : _GEN_7131; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7133 = _GEN_9104 & 4'hd == EntId[3:0] ? dataArray_60_13_cachedata_MPORT_data : _GEN_7132; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7134 = _GEN_9104 & 4'he == EntId[3:0] ? dataArray_60_14_cachedata_MPORT_data : _GEN_7133; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7135 = _GEN_9104 & 4'hf == EntId[3:0] ? dataArray_60_15_cachedata_MPORT_data : _GEN_7134; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7136 = _GEN_9136 & 4'h0 == EntId[3:0] ? dataArray_61_0_cachedata_MPORT_data : _GEN_7135; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7137 = _GEN_9136 & 4'h1 == EntId[3:0] ? dataArray_61_1_cachedata_MPORT_data : _GEN_7136; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7138 = _GEN_9136 & 4'h2 == EntId[3:0] ? dataArray_61_2_cachedata_MPORT_data : _GEN_7137; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7139 = _GEN_9136 & 4'h3 == EntId[3:0] ? dataArray_61_3_cachedata_MPORT_data : _GEN_7138; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7140 = _GEN_9136 & 4'h4 == EntId[3:0] ? dataArray_61_4_cachedata_MPORT_data : _GEN_7139; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7141 = _GEN_9136 & 4'h5 == EntId[3:0] ? dataArray_61_5_cachedata_MPORT_data : _GEN_7140; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7142 = _GEN_9136 & 4'h6 == EntId[3:0] ? dataArray_61_6_cachedata_MPORT_data : _GEN_7141; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7143 = _GEN_9136 & 4'h7 == EntId[3:0] ? dataArray_61_7_cachedata_MPORT_data : _GEN_7142; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7144 = _GEN_9136 & 4'h8 == EntId[3:0] ? dataArray_61_8_cachedata_MPORT_data : _GEN_7143; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7145 = _GEN_9136 & 4'h9 == EntId[3:0] ? dataArray_61_9_cachedata_MPORT_data : _GEN_7144; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7146 = _GEN_9136 & 4'ha == EntId[3:0] ? dataArray_61_10_cachedata_MPORT_data : _GEN_7145; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7147 = _GEN_9136 & 4'hb == EntId[3:0] ? dataArray_61_11_cachedata_MPORT_data : _GEN_7146; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7148 = _GEN_9136 & 4'hc == EntId[3:0] ? dataArray_61_12_cachedata_MPORT_data : _GEN_7147; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7149 = _GEN_9136 & 4'hd == EntId[3:0] ? dataArray_61_13_cachedata_MPORT_data : _GEN_7148; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7150 = _GEN_9136 & 4'he == EntId[3:0] ? dataArray_61_14_cachedata_MPORT_data : _GEN_7149; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7151 = _GEN_9136 & 4'hf == EntId[3:0] ? dataArray_61_15_cachedata_MPORT_data : _GEN_7150; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7152 = _GEN_9168 & 4'h0 == EntId[3:0] ? dataArray_62_0_cachedata_MPORT_data : _GEN_7151; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7153 = _GEN_9168 & 4'h1 == EntId[3:0] ? dataArray_62_1_cachedata_MPORT_data : _GEN_7152; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7154 = _GEN_9168 & 4'h2 == EntId[3:0] ? dataArray_62_2_cachedata_MPORT_data : _GEN_7153; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7155 = _GEN_9168 & 4'h3 == EntId[3:0] ? dataArray_62_3_cachedata_MPORT_data : _GEN_7154; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7156 = _GEN_9168 & 4'h4 == EntId[3:0] ? dataArray_62_4_cachedata_MPORT_data : _GEN_7155; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7157 = _GEN_9168 & 4'h5 == EntId[3:0] ? dataArray_62_5_cachedata_MPORT_data : _GEN_7156; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7158 = _GEN_9168 & 4'h6 == EntId[3:0] ? dataArray_62_6_cachedata_MPORT_data : _GEN_7157; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7159 = _GEN_9168 & 4'h7 == EntId[3:0] ? dataArray_62_7_cachedata_MPORT_data : _GEN_7158; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7160 = _GEN_9168 & 4'h8 == EntId[3:0] ? dataArray_62_8_cachedata_MPORT_data : _GEN_7159; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7161 = _GEN_9168 & 4'h9 == EntId[3:0] ? dataArray_62_9_cachedata_MPORT_data : _GEN_7160; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7162 = _GEN_9168 & 4'ha == EntId[3:0] ? dataArray_62_10_cachedata_MPORT_data : _GEN_7161; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7163 = _GEN_9168 & 4'hb == EntId[3:0] ? dataArray_62_11_cachedata_MPORT_data : _GEN_7162; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7164 = _GEN_9168 & 4'hc == EntId[3:0] ? dataArray_62_12_cachedata_MPORT_data : _GEN_7163; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7165 = _GEN_9168 & 4'hd == EntId[3:0] ? dataArray_62_13_cachedata_MPORT_data : _GEN_7164; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7166 = _GEN_9168 & 4'he == EntId[3:0] ? dataArray_62_14_cachedata_MPORT_data : _GEN_7165; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7167 = _GEN_9168 & 4'hf == EntId[3:0] ? dataArray_62_15_cachedata_MPORT_data : _GEN_7166; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7168 = _GEN_9200 & 4'h0 == EntId[3:0] ? dataArray_63_0_cachedata_MPORT_data : _GEN_7167; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7169 = _GEN_9200 & 4'h1 == EntId[3:0] ? dataArray_63_1_cachedata_MPORT_data : _GEN_7168; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7170 = _GEN_9200 & 4'h2 == EntId[3:0] ? dataArray_63_2_cachedata_MPORT_data : _GEN_7169; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7171 = _GEN_9200 & 4'h3 == EntId[3:0] ? dataArray_63_3_cachedata_MPORT_data : _GEN_7170; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7172 = _GEN_9200 & 4'h4 == EntId[3:0] ? dataArray_63_4_cachedata_MPORT_data : _GEN_7171; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7173 = _GEN_9200 & 4'h5 == EntId[3:0] ? dataArray_63_5_cachedata_MPORT_data : _GEN_7172; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7174 = _GEN_9200 & 4'h6 == EntId[3:0] ? dataArray_63_6_cachedata_MPORT_data : _GEN_7173; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7175 = _GEN_9200 & 4'h7 == EntId[3:0] ? dataArray_63_7_cachedata_MPORT_data : _GEN_7174; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7176 = _GEN_9200 & 4'h8 == EntId[3:0] ? dataArray_63_8_cachedata_MPORT_data : _GEN_7175; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7177 = _GEN_9200 & 4'h9 == EntId[3:0] ? dataArray_63_9_cachedata_MPORT_data : _GEN_7176; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7178 = _GEN_9200 & 4'ha == EntId[3:0] ? dataArray_63_10_cachedata_MPORT_data : _GEN_7177; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7179 = _GEN_9200 & 4'hb == EntId[3:0] ? dataArray_63_11_cachedata_MPORT_data : _GEN_7178; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7180 = _GEN_9200 & 4'hc == EntId[3:0] ? dataArray_63_12_cachedata_MPORT_data : _GEN_7179; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7181 = _GEN_9200 & 4'hd == EntId[3:0] ? dataArray_63_13_cachedata_MPORT_data : _GEN_7180; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7182 = _GEN_9200 & 4'he == EntId[3:0] ? dataArray_63_14_cachedata_MPORT_data : _GEN_7181; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_7183 = _GEN_9200 & 4'hf == EntId[3:0] ? dataArray_63_15_cachedata_MPORT_data : _GEN_7182; // @[cache.scala 108:{28,28}]
  assign dataArray_0_0_cachedata_MPORT_en = dataArray_0_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_0_cachedata_MPORT_addr = dataArray_0_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_0_cachedata_MPORT_data = dataArray_0_0[dataArray_0_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_0_MPORT_addr = replace_set;
  assign dataArray_0_0_MPORT_mask = _GEN_7184 & _GEN_7185;
  assign dataArray_0_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_1_cachedata_MPORT_en = dataArray_0_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_1_cachedata_MPORT_addr = dataArray_0_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_1_cachedata_MPORT_data = dataArray_0_1[dataArray_0_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_1_MPORT_addr = replace_set;
  assign dataArray_0_1_MPORT_mask = _GEN_7184 & _GEN_7187;
  assign dataArray_0_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_2_cachedata_MPORT_en = dataArray_0_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_2_cachedata_MPORT_addr = dataArray_0_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_2_cachedata_MPORT_data = dataArray_0_2[dataArray_0_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_2_MPORT_addr = replace_set;
  assign dataArray_0_2_MPORT_mask = _GEN_7184 & _GEN_7189;
  assign dataArray_0_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_3_cachedata_MPORT_en = dataArray_0_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_3_cachedata_MPORT_addr = dataArray_0_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_3_cachedata_MPORT_data = dataArray_0_3[dataArray_0_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_3_MPORT_addr = replace_set;
  assign dataArray_0_3_MPORT_mask = _GEN_7184 & _GEN_7191;
  assign dataArray_0_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_4_cachedata_MPORT_en = dataArray_0_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_4_cachedata_MPORT_addr = dataArray_0_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_4_cachedata_MPORT_data = dataArray_0_4[dataArray_0_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_4_MPORT_addr = replace_set;
  assign dataArray_0_4_MPORT_mask = _GEN_7184 & _GEN_7193;
  assign dataArray_0_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_5_cachedata_MPORT_en = dataArray_0_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_5_cachedata_MPORT_addr = dataArray_0_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_5_cachedata_MPORT_data = dataArray_0_5[dataArray_0_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_5_MPORT_addr = replace_set;
  assign dataArray_0_5_MPORT_mask = _GEN_7184 & _GEN_7195;
  assign dataArray_0_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_6_cachedata_MPORT_en = dataArray_0_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_6_cachedata_MPORT_addr = dataArray_0_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_6_cachedata_MPORT_data = dataArray_0_6[dataArray_0_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_6_MPORT_addr = replace_set;
  assign dataArray_0_6_MPORT_mask = _GEN_7184 & _GEN_7197;
  assign dataArray_0_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_7_cachedata_MPORT_en = dataArray_0_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_7_cachedata_MPORT_addr = dataArray_0_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_7_cachedata_MPORT_data = dataArray_0_7[dataArray_0_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_7_MPORT_addr = replace_set;
  assign dataArray_0_7_MPORT_mask = _GEN_7184 & _GEN_7199;
  assign dataArray_0_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_8_cachedata_MPORT_en = dataArray_0_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_8_cachedata_MPORT_addr = dataArray_0_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_8_cachedata_MPORT_data = dataArray_0_8[dataArray_0_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_8_MPORT_addr = replace_set;
  assign dataArray_0_8_MPORT_mask = _GEN_7184 & _GEN_7201;
  assign dataArray_0_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_9_cachedata_MPORT_en = dataArray_0_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_9_cachedata_MPORT_addr = dataArray_0_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_9_cachedata_MPORT_data = dataArray_0_9[dataArray_0_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_9_MPORT_addr = replace_set;
  assign dataArray_0_9_MPORT_mask = _GEN_7184 & _GEN_7203;
  assign dataArray_0_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_10_cachedata_MPORT_en = dataArray_0_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_10_cachedata_MPORT_addr = dataArray_0_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_10_cachedata_MPORT_data = dataArray_0_10[dataArray_0_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_10_MPORT_addr = replace_set;
  assign dataArray_0_10_MPORT_mask = _GEN_7184 & _GEN_7205;
  assign dataArray_0_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_11_cachedata_MPORT_en = dataArray_0_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_11_cachedata_MPORT_addr = dataArray_0_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_11_cachedata_MPORT_data = dataArray_0_11[dataArray_0_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_11_MPORT_addr = replace_set;
  assign dataArray_0_11_MPORT_mask = _GEN_7184 & _GEN_7207;
  assign dataArray_0_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_12_cachedata_MPORT_en = dataArray_0_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_12_cachedata_MPORT_addr = dataArray_0_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_12_cachedata_MPORT_data = dataArray_0_12[dataArray_0_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_12_MPORT_addr = replace_set;
  assign dataArray_0_12_MPORT_mask = _GEN_7184 & _GEN_7209;
  assign dataArray_0_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_13_cachedata_MPORT_en = dataArray_0_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_13_cachedata_MPORT_addr = dataArray_0_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_13_cachedata_MPORT_data = dataArray_0_13[dataArray_0_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_13_MPORT_addr = replace_set;
  assign dataArray_0_13_MPORT_mask = _GEN_7184 & _GEN_7211;
  assign dataArray_0_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_14_cachedata_MPORT_en = dataArray_0_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_14_cachedata_MPORT_addr = dataArray_0_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_14_cachedata_MPORT_data = dataArray_0_14[dataArray_0_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_14_MPORT_addr = replace_set;
  assign dataArray_0_14_MPORT_mask = _GEN_7184 & _GEN_7213;
  assign dataArray_0_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_15_cachedata_MPORT_en = dataArray_0_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_15_cachedata_MPORT_addr = dataArray_0_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_15_cachedata_MPORT_data = dataArray_0_15[dataArray_0_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_15_MPORT_addr = replace_set;
  assign dataArray_0_15_MPORT_mask = _GEN_7184 & _GEN_7215;
  assign dataArray_0_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_0_cachedata_MPORT_en = dataArray_1_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_0_cachedata_MPORT_addr = dataArray_1_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_0_cachedata_MPORT_data = dataArray_1_0[dataArray_1_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_0_MPORT_addr = replace_set;
  assign dataArray_1_0_MPORT_mask = _GEN_7216 & _GEN_7185;
  assign dataArray_1_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_1_cachedata_MPORT_en = dataArray_1_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_1_cachedata_MPORT_addr = dataArray_1_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_1_cachedata_MPORT_data = dataArray_1_1[dataArray_1_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_1_MPORT_addr = replace_set;
  assign dataArray_1_1_MPORT_mask = _GEN_7216 & _GEN_7187;
  assign dataArray_1_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_2_cachedata_MPORT_en = dataArray_1_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_2_cachedata_MPORT_addr = dataArray_1_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_2_cachedata_MPORT_data = dataArray_1_2[dataArray_1_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_2_MPORT_addr = replace_set;
  assign dataArray_1_2_MPORT_mask = _GEN_7216 & _GEN_7189;
  assign dataArray_1_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_3_cachedata_MPORT_en = dataArray_1_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_3_cachedata_MPORT_addr = dataArray_1_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_3_cachedata_MPORT_data = dataArray_1_3[dataArray_1_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_3_MPORT_addr = replace_set;
  assign dataArray_1_3_MPORT_mask = _GEN_7216 & _GEN_7191;
  assign dataArray_1_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_4_cachedata_MPORT_en = dataArray_1_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_4_cachedata_MPORT_addr = dataArray_1_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_4_cachedata_MPORT_data = dataArray_1_4[dataArray_1_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_4_MPORT_addr = replace_set;
  assign dataArray_1_4_MPORT_mask = _GEN_7216 & _GEN_7193;
  assign dataArray_1_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_5_cachedata_MPORT_en = dataArray_1_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_5_cachedata_MPORT_addr = dataArray_1_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_5_cachedata_MPORT_data = dataArray_1_5[dataArray_1_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_5_MPORT_addr = replace_set;
  assign dataArray_1_5_MPORT_mask = _GEN_7216 & _GEN_7195;
  assign dataArray_1_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_6_cachedata_MPORT_en = dataArray_1_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_6_cachedata_MPORT_addr = dataArray_1_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_6_cachedata_MPORT_data = dataArray_1_6[dataArray_1_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_6_MPORT_addr = replace_set;
  assign dataArray_1_6_MPORT_mask = _GEN_7216 & _GEN_7197;
  assign dataArray_1_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_7_cachedata_MPORT_en = dataArray_1_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_7_cachedata_MPORT_addr = dataArray_1_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_7_cachedata_MPORT_data = dataArray_1_7[dataArray_1_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_7_MPORT_addr = replace_set;
  assign dataArray_1_7_MPORT_mask = _GEN_7216 & _GEN_7199;
  assign dataArray_1_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_8_cachedata_MPORT_en = dataArray_1_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_8_cachedata_MPORT_addr = dataArray_1_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_8_cachedata_MPORT_data = dataArray_1_8[dataArray_1_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_8_MPORT_addr = replace_set;
  assign dataArray_1_8_MPORT_mask = _GEN_7216 & _GEN_7201;
  assign dataArray_1_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_9_cachedata_MPORT_en = dataArray_1_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_9_cachedata_MPORT_addr = dataArray_1_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_9_cachedata_MPORT_data = dataArray_1_9[dataArray_1_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_9_MPORT_addr = replace_set;
  assign dataArray_1_9_MPORT_mask = _GEN_7216 & _GEN_7203;
  assign dataArray_1_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_10_cachedata_MPORT_en = dataArray_1_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_10_cachedata_MPORT_addr = dataArray_1_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_10_cachedata_MPORT_data = dataArray_1_10[dataArray_1_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_10_MPORT_addr = replace_set;
  assign dataArray_1_10_MPORT_mask = _GEN_7216 & _GEN_7205;
  assign dataArray_1_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_11_cachedata_MPORT_en = dataArray_1_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_11_cachedata_MPORT_addr = dataArray_1_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_11_cachedata_MPORT_data = dataArray_1_11[dataArray_1_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_11_MPORT_addr = replace_set;
  assign dataArray_1_11_MPORT_mask = _GEN_7216 & _GEN_7207;
  assign dataArray_1_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_12_cachedata_MPORT_en = dataArray_1_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_12_cachedata_MPORT_addr = dataArray_1_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_12_cachedata_MPORT_data = dataArray_1_12[dataArray_1_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_12_MPORT_addr = replace_set;
  assign dataArray_1_12_MPORT_mask = _GEN_7216 & _GEN_7209;
  assign dataArray_1_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_13_cachedata_MPORT_en = dataArray_1_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_13_cachedata_MPORT_addr = dataArray_1_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_13_cachedata_MPORT_data = dataArray_1_13[dataArray_1_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_13_MPORT_addr = replace_set;
  assign dataArray_1_13_MPORT_mask = _GEN_7216 & _GEN_7211;
  assign dataArray_1_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_14_cachedata_MPORT_en = dataArray_1_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_14_cachedata_MPORT_addr = dataArray_1_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_14_cachedata_MPORT_data = dataArray_1_14[dataArray_1_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_14_MPORT_addr = replace_set;
  assign dataArray_1_14_MPORT_mask = _GEN_7216 & _GEN_7213;
  assign dataArray_1_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_15_cachedata_MPORT_en = dataArray_1_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_15_cachedata_MPORT_addr = dataArray_1_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_15_cachedata_MPORT_data = dataArray_1_15[dataArray_1_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_15_MPORT_addr = replace_set;
  assign dataArray_1_15_MPORT_mask = _GEN_7216 & _GEN_7215;
  assign dataArray_1_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_0_cachedata_MPORT_en = dataArray_2_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_0_cachedata_MPORT_addr = dataArray_2_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_0_cachedata_MPORT_data = dataArray_2_0[dataArray_2_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_0_MPORT_addr = replace_set;
  assign dataArray_2_0_MPORT_mask = _GEN_7248 & _GEN_7185;
  assign dataArray_2_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_1_cachedata_MPORT_en = dataArray_2_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_1_cachedata_MPORT_addr = dataArray_2_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_1_cachedata_MPORT_data = dataArray_2_1[dataArray_2_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_1_MPORT_addr = replace_set;
  assign dataArray_2_1_MPORT_mask = _GEN_7248 & _GEN_7187;
  assign dataArray_2_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_2_cachedata_MPORT_en = dataArray_2_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_2_cachedata_MPORT_addr = dataArray_2_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_2_cachedata_MPORT_data = dataArray_2_2[dataArray_2_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_2_MPORT_addr = replace_set;
  assign dataArray_2_2_MPORT_mask = _GEN_7248 & _GEN_7189;
  assign dataArray_2_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_3_cachedata_MPORT_en = dataArray_2_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_3_cachedata_MPORT_addr = dataArray_2_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_3_cachedata_MPORT_data = dataArray_2_3[dataArray_2_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_3_MPORT_addr = replace_set;
  assign dataArray_2_3_MPORT_mask = _GEN_7248 & _GEN_7191;
  assign dataArray_2_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_4_cachedata_MPORT_en = dataArray_2_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_4_cachedata_MPORT_addr = dataArray_2_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_4_cachedata_MPORT_data = dataArray_2_4[dataArray_2_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_4_MPORT_addr = replace_set;
  assign dataArray_2_4_MPORT_mask = _GEN_7248 & _GEN_7193;
  assign dataArray_2_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_5_cachedata_MPORT_en = dataArray_2_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_5_cachedata_MPORT_addr = dataArray_2_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_5_cachedata_MPORT_data = dataArray_2_5[dataArray_2_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_5_MPORT_addr = replace_set;
  assign dataArray_2_5_MPORT_mask = _GEN_7248 & _GEN_7195;
  assign dataArray_2_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_6_cachedata_MPORT_en = dataArray_2_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_6_cachedata_MPORT_addr = dataArray_2_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_6_cachedata_MPORT_data = dataArray_2_6[dataArray_2_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_6_MPORT_addr = replace_set;
  assign dataArray_2_6_MPORT_mask = _GEN_7248 & _GEN_7197;
  assign dataArray_2_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_7_cachedata_MPORT_en = dataArray_2_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_7_cachedata_MPORT_addr = dataArray_2_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_7_cachedata_MPORT_data = dataArray_2_7[dataArray_2_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_7_MPORT_addr = replace_set;
  assign dataArray_2_7_MPORT_mask = _GEN_7248 & _GEN_7199;
  assign dataArray_2_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_8_cachedata_MPORT_en = dataArray_2_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_8_cachedata_MPORT_addr = dataArray_2_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_8_cachedata_MPORT_data = dataArray_2_8[dataArray_2_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_8_MPORT_addr = replace_set;
  assign dataArray_2_8_MPORT_mask = _GEN_7248 & _GEN_7201;
  assign dataArray_2_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_9_cachedata_MPORT_en = dataArray_2_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_9_cachedata_MPORT_addr = dataArray_2_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_9_cachedata_MPORT_data = dataArray_2_9[dataArray_2_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_9_MPORT_addr = replace_set;
  assign dataArray_2_9_MPORT_mask = _GEN_7248 & _GEN_7203;
  assign dataArray_2_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_10_cachedata_MPORT_en = dataArray_2_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_10_cachedata_MPORT_addr = dataArray_2_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_10_cachedata_MPORT_data = dataArray_2_10[dataArray_2_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_10_MPORT_addr = replace_set;
  assign dataArray_2_10_MPORT_mask = _GEN_7248 & _GEN_7205;
  assign dataArray_2_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_11_cachedata_MPORT_en = dataArray_2_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_11_cachedata_MPORT_addr = dataArray_2_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_11_cachedata_MPORT_data = dataArray_2_11[dataArray_2_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_11_MPORT_addr = replace_set;
  assign dataArray_2_11_MPORT_mask = _GEN_7248 & _GEN_7207;
  assign dataArray_2_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_12_cachedata_MPORT_en = dataArray_2_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_12_cachedata_MPORT_addr = dataArray_2_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_12_cachedata_MPORT_data = dataArray_2_12[dataArray_2_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_12_MPORT_addr = replace_set;
  assign dataArray_2_12_MPORT_mask = _GEN_7248 & _GEN_7209;
  assign dataArray_2_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_13_cachedata_MPORT_en = dataArray_2_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_13_cachedata_MPORT_addr = dataArray_2_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_13_cachedata_MPORT_data = dataArray_2_13[dataArray_2_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_13_MPORT_addr = replace_set;
  assign dataArray_2_13_MPORT_mask = _GEN_7248 & _GEN_7211;
  assign dataArray_2_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_14_cachedata_MPORT_en = dataArray_2_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_14_cachedata_MPORT_addr = dataArray_2_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_14_cachedata_MPORT_data = dataArray_2_14[dataArray_2_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_14_MPORT_addr = replace_set;
  assign dataArray_2_14_MPORT_mask = _GEN_7248 & _GEN_7213;
  assign dataArray_2_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_15_cachedata_MPORT_en = dataArray_2_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_15_cachedata_MPORT_addr = dataArray_2_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_15_cachedata_MPORT_data = dataArray_2_15[dataArray_2_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_15_MPORT_addr = replace_set;
  assign dataArray_2_15_MPORT_mask = _GEN_7248 & _GEN_7215;
  assign dataArray_2_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_0_cachedata_MPORT_en = dataArray_3_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_0_cachedata_MPORT_addr = dataArray_3_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_0_cachedata_MPORT_data = dataArray_3_0[dataArray_3_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_0_MPORT_addr = replace_set;
  assign dataArray_3_0_MPORT_mask = _GEN_7280 & _GEN_7185;
  assign dataArray_3_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_1_cachedata_MPORT_en = dataArray_3_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_1_cachedata_MPORT_addr = dataArray_3_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_1_cachedata_MPORT_data = dataArray_3_1[dataArray_3_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_1_MPORT_addr = replace_set;
  assign dataArray_3_1_MPORT_mask = _GEN_7280 & _GEN_7187;
  assign dataArray_3_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_2_cachedata_MPORT_en = dataArray_3_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_2_cachedata_MPORT_addr = dataArray_3_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_2_cachedata_MPORT_data = dataArray_3_2[dataArray_3_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_2_MPORT_addr = replace_set;
  assign dataArray_3_2_MPORT_mask = _GEN_7280 & _GEN_7189;
  assign dataArray_3_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_3_cachedata_MPORT_en = dataArray_3_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_3_cachedata_MPORT_addr = dataArray_3_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_3_cachedata_MPORT_data = dataArray_3_3[dataArray_3_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_3_MPORT_addr = replace_set;
  assign dataArray_3_3_MPORT_mask = _GEN_7280 & _GEN_7191;
  assign dataArray_3_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_4_cachedata_MPORT_en = dataArray_3_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_4_cachedata_MPORT_addr = dataArray_3_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_4_cachedata_MPORT_data = dataArray_3_4[dataArray_3_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_4_MPORT_addr = replace_set;
  assign dataArray_3_4_MPORT_mask = _GEN_7280 & _GEN_7193;
  assign dataArray_3_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_5_cachedata_MPORT_en = dataArray_3_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_5_cachedata_MPORT_addr = dataArray_3_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_5_cachedata_MPORT_data = dataArray_3_5[dataArray_3_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_5_MPORT_addr = replace_set;
  assign dataArray_3_5_MPORT_mask = _GEN_7280 & _GEN_7195;
  assign dataArray_3_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_6_cachedata_MPORT_en = dataArray_3_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_6_cachedata_MPORT_addr = dataArray_3_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_6_cachedata_MPORT_data = dataArray_3_6[dataArray_3_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_6_MPORT_addr = replace_set;
  assign dataArray_3_6_MPORT_mask = _GEN_7280 & _GEN_7197;
  assign dataArray_3_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_7_cachedata_MPORT_en = dataArray_3_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_7_cachedata_MPORT_addr = dataArray_3_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_7_cachedata_MPORT_data = dataArray_3_7[dataArray_3_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_7_MPORT_addr = replace_set;
  assign dataArray_3_7_MPORT_mask = _GEN_7280 & _GEN_7199;
  assign dataArray_3_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_8_cachedata_MPORT_en = dataArray_3_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_8_cachedata_MPORT_addr = dataArray_3_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_8_cachedata_MPORT_data = dataArray_3_8[dataArray_3_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_8_MPORT_addr = replace_set;
  assign dataArray_3_8_MPORT_mask = _GEN_7280 & _GEN_7201;
  assign dataArray_3_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_9_cachedata_MPORT_en = dataArray_3_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_9_cachedata_MPORT_addr = dataArray_3_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_9_cachedata_MPORT_data = dataArray_3_9[dataArray_3_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_9_MPORT_addr = replace_set;
  assign dataArray_3_9_MPORT_mask = _GEN_7280 & _GEN_7203;
  assign dataArray_3_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_10_cachedata_MPORT_en = dataArray_3_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_10_cachedata_MPORT_addr = dataArray_3_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_10_cachedata_MPORT_data = dataArray_3_10[dataArray_3_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_10_MPORT_addr = replace_set;
  assign dataArray_3_10_MPORT_mask = _GEN_7280 & _GEN_7205;
  assign dataArray_3_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_11_cachedata_MPORT_en = dataArray_3_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_11_cachedata_MPORT_addr = dataArray_3_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_11_cachedata_MPORT_data = dataArray_3_11[dataArray_3_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_11_MPORT_addr = replace_set;
  assign dataArray_3_11_MPORT_mask = _GEN_7280 & _GEN_7207;
  assign dataArray_3_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_12_cachedata_MPORT_en = dataArray_3_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_12_cachedata_MPORT_addr = dataArray_3_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_12_cachedata_MPORT_data = dataArray_3_12[dataArray_3_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_12_MPORT_addr = replace_set;
  assign dataArray_3_12_MPORT_mask = _GEN_7280 & _GEN_7209;
  assign dataArray_3_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_13_cachedata_MPORT_en = dataArray_3_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_13_cachedata_MPORT_addr = dataArray_3_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_13_cachedata_MPORT_data = dataArray_3_13[dataArray_3_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_13_MPORT_addr = replace_set;
  assign dataArray_3_13_MPORT_mask = _GEN_7280 & _GEN_7211;
  assign dataArray_3_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_14_cachedata_MPORT_en = dataArray_3_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_14_cachedata_MPORT_addr = dataArray_3_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_14_cachedata_MPORT_data = dataArray_3_14[dataArray_3_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_14_MPORT_addr = replace_set;
  assign dataArray_3_14_MPORT_mask = _GEN_7280 & _GEN_7213;
  assign dataArray_3_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_15_cachedata_MPORT_en = dataArray_3_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_15_cachedata_MPORT_addr = dataArray_3_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_15_cachedata_MPORT_data = dataArray_3_15[dataArray_3_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_15_MPORT_addr = replace_set;
  assign dataArray_3_15_MPORT_mask = _GEN_7280 & _GEN_7215;
  assign dataArray_3_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_0_cachedata_MPORT_en = dataArray_4_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_0_cachedata_MPORT_addr = dataArray_4_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_0_cachedata_MPORT_data = dataArray_4_0[dataArray_4_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_0_MPORT_addr = replace_set;
  assign dataArray_4_0_MPORT_mask = _GEN_7312 & _GEN_7185;
  assign dataArray_4_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_1_cachedata_MPORT_en = dataArray_4_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_1_cachedata_MPORT_addr = dataArray_4_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_1_cachedata_MPORT_data = dataArray_4_1[dataArray_4_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_1_MPORT_addr = replace_set;
  assign dataArray_4_1_MPORT_mask = _GEN_7312 & _GEN_7187;
  assign dataArray_4_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_2_cachedata_MPORT_en = dataArray_4_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_2_cachedata_MPORT_addr = dataArray_4_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_2_cachedata_MPORT_data = dataArray_4_2[dataArray_4_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_2_MPORT_addr = replace_set;
  assign dataArray_4_2_MPORT_mask = _GEN_7312 & _GEN_7189;
  assign dataArray_4_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_3_cachedata_MPORT_en = dataArray_4_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_3_cachedata_MPORT_addr = dataArray_4_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_3_cachedata_MPORT_data = dataArray_4_3[dataArray_4_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_3_MPORT_addr = replace_set;
  assign dataArray_4_3_MPORT_mask = _GEN_7312 & _GEN_7191;
  assign dataArray_4_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_4_cachedata_MPORT_en = dataArray_4_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_4_cachedata_MPORT_addr = dataArray_4_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_4_cachedata_MPORT_data = dataArray_4_4[dataArray_4_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_4_MPORT_addr = replace_set;
  assign dataArray_4_4_MPORT_mask = _GEN_7312 & _GEN_7193;
  assign dataArray_4_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_5_cachedata_MPORT_en = dataArray_4_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_5_cachedata_MPORT_addr = dataArray_4_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_5_cachedata_MPORT_data = dataArray_4_5[dataArray_4_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_5_MPORT_addr = replace_set;
  assign dataArray_4_5_MPORT_mask = _GEN_7312 & _GEN_7195;
  assign dataArray_4_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_6_cachedata_MPORT_en = dataArray_4_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_6_cachedata_MPORT_addr = dataArray_4_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_6_cachedata_MPORT_data = dataArray_4_6[dataArray_4_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_6_MPORT_addr = replace_set;
  assign dataArray_4_6_MPORT_mask = _GEN_7312 & _GEN_7197;
  assign dataArray_4_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_7_cachedata_MPORT_en = dataArray_4_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_7_cachedata_MPORT_addr = dataArray_4_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_7_cachedata_MPORT_data = dataArray_4_7[dataArray_4_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_7_MPORT_addr = replace_set;
  assign dataArray_4_7_MPORT_mask = _GEN_7312 & _GEN_7199;
  assign dataArray_4_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_8_cachedata_MPORT_en = dataArray_4_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_8_cachedata_MPORT_addr = dataArray_4_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_8_cachedata_MPORT_data = dataArray_4_8[dataArray_4_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_8_MPORT_addr = replace_set;
  assign dataArray_4_8_MPORT_mask = _GEN_7312 & _GEN_7201;
  assign dataArray_4_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_9_cachedata_MPORT_en = dataArray_4_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_9_cachedata_MPORT_addr = dataArray_4_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_9_cachedata_MPORT_data = dataArray_4_9[dataArray_4_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_9_MPORT_addr = replace_set;
  assign dataArray_4_9_MPORT_mask = _GEN_7312 & _GEN_7203;
  assign dataArray_4_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_10_cachedata_MPORT_en = dataArray_4_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_10_cachedata_MPORT_addr = dataArray_4_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_10_cachedata_MPORT_data = dataArray_4_10[dataArray_4_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_10_MPORT_addr = replace_set;
  assign dataArray_4_10_MPORT_mask = _GEN_7312 & _GEN_7205;
  assign dataArray_4_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_11_cachedata_MPORT_en = dataArray_4_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_11_cachedata_MPORT_addr = dataArray_4_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_11_cachedata_MPORT_data = dataArray_4_11[dataArray_4_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_11_MPORT_addr = replace_set;
  assign dataArray_4_11_MPORT_mask = _GEN_7312 & _GEN_7207;
  assign dataArray_4_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_12_cachedata_MPORT_en = dataArray_4_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_12_cachedata_MPORT_addr = dataArray_4_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_12_cachedata_MPORT_data = dataArray_4_12[dataArray_4_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_12_MPORT_addr = replace_set;
  assign dataArray_4_12_MPORT_mask = _GEN_7312 & _GEN_7209;
  assign dataArray_4_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_13_cachedata_MPORT_en = dataArray_4_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_13_cachedata_MPORT_addr = dataArray_4_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_13_cachedata_MPORT_data = dataArray_4_13[dataArray_4_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_13_MPORT_addr = replace_set;
  assign dataArray_4_13_MPORT_mask = _GEN_7312 & _GEN_7211;
  assign dataArray_4_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_14_cachedata_MPORT_en = dataArray_4_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_14_cachedata_MPORT_addr = dataArray_4_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_14_cachedata_MPORT_data = dataArray_4_14[dataArray_4_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_14_MPORT_addr = replace_set;
  assign dataArray_4_14_MPORT_mask = _GEN_7312 & _GEN_7213;
  assign dataArray_4_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_15_cachedata_MPORT_en = dataArray_4_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_15_cachedata_MPORT_addr = dataArray_4_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_15_cachedata_MPORT_data = dataArray_4_15[dataArray_4_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_15_MPORT_addr = replace_set;
  assign dataArray_4_15_MPORT_mask = _GEN_7312 & _GEN_7215;
  assign dataArray_4_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_0_cachedata_MPORT_en = dataArray_5_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_0_cachedata_MPORT_addr = dataArray_5_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_0_cachedata_MPORT_data = dataArray_5_0[dataArray_5_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_0_MPORT_addr = replace_set;
  assign dataArray_5_0_MPORT_mask = _GEN_7344 & _GEN_7185;
  assign dataArray_5_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_1_cachedata_MPORT_en = dataArray_5_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_1_cachedata_MPORT_addr = dataArray_5_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_1_cachedata_MPORT_data = dataArray_5_1[dataArray_5_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_1_MPORT_addr = replace_set;
  assign dataArray_5_1_MPORT_mask = _GEN_7344 & _GEN_7187;
  assign dataArray_5_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_2_cachedata_MPORT_en = dataArray_5_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_2_cachedata_MPORT_addr = dataArray_5_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_2_cachedata_MPORT_data = dataArray_5_2[dataArray_5_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_2_MPORT_addr = replace_set;
  assign dataArray_5_2_MPORT_mask = _GEN_7344 & _GEN_7189;
  assign dataArray_5_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_3_cachedata_MPORT_en = dataArray_5_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_3_cachedata_MPORT_addr = dataArray_5_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_3_cachedata_MPORT_data = dataArray_5_3[dataArray_5_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_3_MPORT_addr = replace_set;
  assign dataArray_5_3_MPORT_mask = _GEN_7344 & _GEN_7191;
  assign dataArray_5_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_4_cachedata_MPORT_en = dataArray_5_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_4_cachedata_MPORT_addr = dataArray_5_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_4_cachedata_MPORT_data = dataArray_5_4[dataArray_5_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_4_MPORT_addr = replace_set;
  assign dataArray_5_4_MPORT_mask = _GEN_7344 & _GEN_7193;
  assign dataArray_5_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_5_cachedata_MPORT_en = dataArray_5_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_5_cachedata_MPORT_addr = dataArray_5_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_5_cachedata_MPORT_data = dataArray_5_5[dataArray_5_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_5_MPORT_addr = replace_set;
  assign dataArray_5_5_MPORT_mask = _GEN_7344 & _GEN_7195;
  assign dataArray_5_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_6_cachedata_MPORT_en = dataArray_5_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_6_cachedata_MPORT_addr = dataArray_5_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_6_cachedata_MPORT_data = dataArray_5_6[dataArray_5_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_6_MPORT_addr = replace_set;
  assign dataArray_5_6_MPORT_mask = _GEN_7344 & _GEN_7197;
  assign dataArray_5_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_7_cachedata_MPORT_en = dataArray_5_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_7_cachedata_MPORT_addr = dataArray_5_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_7_cachedata_MPORT_data = dataArray_5_7[dataArray_5_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_7_MPORT_addr = replace_set;
  assign dataArray_5_7_MPORT_mask = _GEN_7344 & _GEN_7199;
  assign dataArray_5_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_8_cachedata_MPORT_en = dataArray_5_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_8_cachedata_MPORT_addr = dataArray_5_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_8_cachedata_MPORT_data = dataArray_5_8[dataArray_5_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_8_MPORT_addr = replace_set;
  assign dataArray_5_8_MPORT_mask = _GEN_7344 & _GEN_7201;
  assign dataArray_5_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_9_cachedata_MPORT_en = dataArray_5_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_9_cachedata_MPORT_addr = dataArray_5_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_9_cachedata_MPORT_data = dataArray_5_9[dataArray_5_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_9_MPORT_addr = replace_set;
  assign dataArray_5_9_MPORT_mask = _GEN_7344 & _GEN_7203;
  assign dataArray_5_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_10_cachedata_MPORT_en = dataArray_5_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_10_cachedata_MPORT_addr = dataArray_5_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_10_cachedata_MPORT_data = dataArray_5_10[dataArray_5_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_10_MPORT_addr = replace_set;
  assign dataArray_5_10_MPORT_mask = _GEN_7344 & _GEN_7205;
  assign dataArray_5_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_11_cachedata_MPORT_en = dataArray_5_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_11_cachedata_MPORT_addr = dataArray_5_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_11_cachedata_MPORT_data = dataArray_5_11[dataArray_5_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_11_MPORT_addr = replace_set;
  assign dataArray_5_11_MPORT_mask = _GEN_7344 & _GEN_7207;
  assign dataArray_5_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_12_cachedata_MPORT_en = dataArray_5_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_12_cachedata_MPORT_addr = dataArray_5_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_12_cachedata_MPORT_data = dataArray_5_12[dataArray_5_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_12_MPORT_addr = replace_set;
  assign dataArray_5_12_MPORT_mask = _GEN_7344 & _GEN_7209;
  assign dataArray_5_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_13_cachedata_MPORT_en = dataArray_5_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_13_cachedata_MPORT_addr = dataArray_5_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_13_cachedata_MPORT_data = dataArray_5_13[dataArray_5_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_13_MPORT_addr = replace_set;
  assign dataArray_5_13_MPORT_mask = _GEN_7344 & _GEN_7211;
  assign dataArray_5_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_14_cachedata_MPORT_en = dataArray_5_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_14_cachedata_MPORT_addr = dataArray_5_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_14_cachedata_MPORT_data = dataArray_5_14[dataArray_5_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_14_MPORT_addr = replace_set;
  assign dataArray_5_14_MPORT_mask = _GEN_7344 & _GEN_7213;
  assign dataArray_5_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_15_cachedata_MPORT_en = dataArray_5_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_15_cachedata_MPORT_addr = dataArray_5_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_15_cachedata_MPORT_data = dataArray_5_15[dataArray_5_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_15_MPORT_addr = replace_set;
  assign dataArray_5_15_MPORT_mask = _GEN_7344 & _GEN_7215;
  assign dataArray_5_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_0_cachedata_MPORT_en = dataArray_6_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_0_cachedata_MPORT_addr = dataArray_6_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_0_cachedata_MPORT_data = dataArray_6_0[dataArray_6_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_0_MPORT_addr = replace_set;
  assign dataArray_6_0_MPORT_mask = _GEN_7376 & _GEN_7185;
  assign dataArray_6_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_1_cachedata_MPORT_en = dataArray_6_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_1_cachedata_MPORT_addr = dataArray_6_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_1_cachedata_MPORT_data = dataArray_6_1[dataArray_6_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_1_MPORT_addr = replace_set;
  assign dataArray_6_1_MPORT_mask = _GEN_7376 & _GEN_7187;
  assign dataArray_6_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_2_cachedata_MPORT_en = dataArray_6_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_2_cachedata_MPORT_addr = dataArray_6_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_2_cachedata_MPORT_data = dataArray_6_2[dataArray_6_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_2_MPORT_addr = replace_set;
  assign dataArray_6_2_MPORT_mask = _GEN_7376 & _GEN_7189;
  assign dataArray_6_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_3_cachedata_MPORT_en = dataArray_6_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_3_cachedata_MPORT_addr = dataArray_6_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_3_cachedata_MPORT_data = dataArray_6_3[dataArray_6_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_3_MPORT_addr = replace_set;
  assign dataArray_6_3_MPORT_mask = _GEN_7376 & _GEN_7191;
  assign dataArray_6_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_4_cachedata_MPORT_en = dataArray_6_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_4_cachedata_MPORT_addr = dataArray_6_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_4_cachedata_MPORT_data = dataArray_6_4[dataArray_6_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_4_MPORT_addr = replace_set;
  assign dataArray_6_4_MPORT_mask = _GEN_7376 & _GEN_7193;
  assign dataArray_6_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_5_cachedata_MPORT_en = dataArray_6_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_5_cachedata_MPORT_addr = dataArray_6_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_5_cachedata_MPORT_data = dataArray_6_5[dataArray_6_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_5_MPORT_addr = replace_set;
  assign dataArray_6_5_MPORT_mask = _GEN_7376 & _GEN_7195;
  assign dataArray_6_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_6_cachedata_MPORT_en = dataArray_6_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_6_cachedata_MPORT_addr = dataArray_6_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_6_cachedata_MPORT_data = dataArray_6_6[dataArray_6_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_6_MPORT_addr = replace_set;
  assign dataArray_6_6_MPORT_mask = _GEN_7376 & _GEN_7197;
  assign dataArray_6_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_7_cachedata_MPORT_en = dataArray_6_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_7_cachedata_MPORT_addr = dataArray_6_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_7_cachedata_MPORT_data = dataArray_6_7[dataArray_6_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_7_MPORT_addr = replace_set;
  assign dataArray_6_7_MPORT_mask = _GEN_7376 & _GEN_7199;
  assign dataArray_6_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_8_cachedata_MPORT_en = dataArray_6_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_8_cachedata_MPORT_addr = dataArray_6_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_8_cachedata_MPORT_data = dataArray_6_8[dataArray_6_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_8_MPORT_addr = replace_set;
  assign dataArray_6_8_MPORT_mask = _GEN_7376 & _GEN_7201;
  assign dataArray_6_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_9_cachedata_MPORT_en = dataArray_6_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_9_cachedata_MPORT_addr = dataArray_6_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_9_cachedata_MPORT_data = dataArray_6_9[dataArray_6_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_9_MPORT_addr = replace_set;
  assign dataArray_6_9_MPORT_mask = _GEN_7376 & _GEN_7203;
  assign dataArray_6_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_10_cachedata_MPORT_en = dataArray_6_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_10_cachedata_MPORT_addr = dataArray_6_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_10_cachedata_MPORT_data = dataArray_6_10[dataArray_6_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_10_MPORT_addr = replace_set;
  assign dataArray_6_10_MPORT_mask = _GEN_7376 & _GEN_7205;
  assign dataArray_6_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_11_cachedata_MPORT_en = dataArray_6_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_11_cachedata_MPORT_addr = dataArray_6_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_11_cachedata_MPORT_data = dataArray_6_11[dataArray_6_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_11_MPORT_addr = replace_set;
  assign dataArray_6_11_MPORT_mask = _GEN_7376 & _GEN_7207;
  assign dataArray_6_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_12_cachedata_MPORT_en = dataArray_6_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_12_cachedata_MPORT_addr = dataArray_6_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_12_cachedata_MPORT_data = dataArray_6_12[dataArray_6_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_12_MPORT_addr = replace_set;
  assign dataArray_6_12_MPORT_mask = _GEN_7376 & _GEN_7209;
  assign dataArray_6_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_13_cachedata_MPORT_en = dataArray_6_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_13_cachedata_MPORT_addr = dataArray_6_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_13_cachedata_MPORT_data = dataArray_6_13[dataArray_6_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_13_MPORT_addr = replace_set;
  assign dataArray_6_13_MPORT_mask = _GEN_7376 & _GEN_7211;
  assign dataArray_6_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_14_cachedata_MPORT_en = dataArray_6_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_14_cachedata_MPORT_addr = dataArray_6_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_14_cachedata_MPORT_data = dataArray_6_14[dataArray_6_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_14_MPORT_addr = replace_set;
  assign dataArray_6_14_MPORT_mask = _GEN_7376 & _GEN_7213;
  assign dataArray_6_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_15_cachedata_MPORT_en = dataArray_6_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_15_cachedata_MPORT_addr = dataArray_6_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_15_cachedata_MPORT_data = dataArray_6_15[dataArray_6_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_15_MPORT_addr = replace_set;
  assign dataArray_6_15_MPORT_mask = _GEN_7376 & _GEN_7215;
  assign dataArray_6_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_0_cachedata_MPORT_en = dataArray_7_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_0_cachedata_MPORT_addr = dataArray_7_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_0_cachedata_MPORT_data = dataArray_7_0[dataArray_7_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_0_MPORT_addr = replace_set;
  assign dataArray_7_0_MPORT_mask = _GEN_7408 & _GEN_7185;
  assign dataArray_7_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_1_cachedata_MPORT_en = dataArray_7_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_1_cachedata_MPORT_addr = dataArray_7_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_1_cachedata_MPORT_data = dataArray_7_1[dataArray_7_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_1_MPORT_addr = replace_set;
  assign dataArray_7_1_MPORT_mask = _GEN_7408 & _GEN_7187;
  assign dataArray_7_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_2_cachedata_MPORT_en = dataArray_7_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_2_cachedata_MPORT_addr = dataArray_7_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_2_cachedata_MPORT_data = dataArray_7_2[dataArray_7_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_2_MPORT_addr = replace_set;
  assign dataArray_7_2_MPORT_mask = _GEN_7408 & _GEN_7189;
  assign dataArray_7_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_3_cachedata_MPORT_en = dataArray_7_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_3_cachedata_MPORT_addr = dataArray_7_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_3_cachedata_MPORT_data = dataArray_7_3[dataArray_7_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_3_MPORT_addr = replace_set;
  assign dataArray_7_3_MPORT_mask = _GEN_7408 & _GEN_7191;
  assign dataArray_7_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_4_cachedata_MPORT_en = dataArray_7_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_4_cachedata_MPORT_addr = dataArray_7_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_4_cachedata_MPORT_data = dataArray_7_4[dataArray_7_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_4_MPORT_addr = replace_set;
  assign dataArray_7_4_MPORT_mask = _GEN_7408 & _GEN_7193;
  assign dataArray_7_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_5_cachedata_MPORT_en = dataArray_7_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_5_cachedata_MPORT_addr = dataArray_7_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_5_cachedata_MPORT_data = dataArray_7_5[dataArray_7_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_5_MPORT_addr = replace_set;
  assign dataArray_7_5_MPORT_mask = _GEN_7408 & _GEN_7195;
  assign dataArray_7_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_6_cachedata_MPORT_en = dataArray_7_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_6_cachedata_MPORT_addr = dataArray_7_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_6_cachedata_MPORT_data = dataArray_7_6[dataArray_7_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_6_MPORT_addr = replace_set;
  assign dataArray_7_6_MPORT_mask = _GEN_7408 & _GEN_7197;
  assign dataArray_7_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_7_cachedata_MPORT_en = dataArray_7_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_7_cachedata_MPORT_addr = dataArray_7_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_7_cachedata_MPORT_data = dataArray_7_7[dataArray_7_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_7_MPORT_addr = replace_set;
  assign dataArray_7_7_MPORT_mask = _GEN_7408 & _GEN_7199;
  assign dataArray_7_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_8_cachedata_MPORT_en = dataArray_7_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_8_cachedata_MPORT_addr = dataArray_7_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_8_cachedata_MPORT_data = dataArray_7_8[dataArray_7_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_8_MPORT_addr = replace_set;
  assign dataArray_7_8_MPORT_mask = _GEN_7408 & _GEN_7201;
  assign dataArray_7_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_9_cachedata_MPORT_en = dataArray_7_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_9_cachedata_MPORT_addr = dataArray_7_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_9_cachedata_MPORT_data = dataArray_7_9[dataArray_7_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_9_MPORT_addr = replace_set;
  assign dataArray_7_9_MPORT_mask = _GEN_7408 & _GEN_7203;
  assign dataArray_7_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_10_cachedata_MPORT_en = dataArray_7_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_10_cachedata_MPORT_addr = dataArray_7_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_10_cachedata_MPORT_data = dataArray_7_10[dataArray_7_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_10_MPORT_addr = replace_set;
  assign dataArray_7_10_MPORT_mask = _GEN_7408 & _GEN_7205;
  assign dataArray_7_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_11_cachedata_MPORT_en = dataArray_7_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_11_cachedata_MPORT_addr = dataArray_7_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_11_cachedata_MPORT_data = dataArray_7_11[dataArray_7_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_11_MPORT_addr = replace_set;
  assign dataArray_7_11_MPORT_mask = _GEN_7408 & _GEN_7207;
  assign dataArray_7_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_12_cachedata_MPORT_en = dataArray_7_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_12_cachedata_MPORT_addr = dataArray_7_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_12_cachedata_MPORT_data = dataArray_7_12[dataArray_7_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_12_MPORT_addr = replace_set;
  assign dataArray_7_12_MPORT_mask = _GEN_7408 & _GEN_7209;
  assign dataArray_7_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_13_cachedata_MPORT_en = dataArray_7_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_13_cachedata_MPORT_addr = dataArray_7_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_13_cachedata_MPORT_data = dataArray_7_13[dataArray_7_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_13_MPORT_addr = replace_set;
  assign dataArray_7_13_MPORT_mask = _GEN_7408 & _GEN_7211;
  assign dataArray_7_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_14_cachedata_MPORT_en = dataArray_7_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_14_cachedata_MPORT_addr = dataArray_7_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_14_cachedata_MPORT_data = dataArray_7_14[dataArray_7_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_14_MPORT_addr = replace_set;
  assign dataArray_7_14_MPORT_mask = _GEN_7408 & _GEN_7213;
  assign dataArray_7_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_15_cachedata_MPORT_en = dataArray_7_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_15_cachedata_MPORT_addr = dataArray_7_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_15_cachedata_MPORT_data = dataArray_7_15[dataArray_7_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_15_MPORT_addr = replace_set;
  assign dataArray_7_15_MPORT_mask = _GEN_7408 & _GEN_7215;
  assign dataArray_7_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_0_cachedata_MPORT_en = dataArray_8_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_0_cachedata_MPORT_addr = dataArray_8_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_0_cachedata_MPORT_data = dataArray_8_0[dataArray_8_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_0_MPORT_addr = replace_set;
  assign dataArray_8_0_MPORT_mask = _GEN_7440 & _GEN_7185;
  assign dataArray_8_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_1_cachedata_MPORT_en = dataArray_8_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_1_cachedata_MPORT_addr = dataArray_8_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_1_cachedata_MPORT_data = dataArray_8_1[dataArray_8_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_1_MPORT_addr = replace_set;
  assign dataArray_8_1_MPORT_mask = _GEN_7440 & _GEN_7187;
  assign dataArray_8_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_2_cachedata_MPORT_en = dataArray_8_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_2_cachedata_MPORT_addr = dataArray_8_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_2_cachedata_MPORT_data = dataArray_8_2[dataArray_8_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_2_MPORT_addr = replace_set;
  assign dataArray_8_2_MPORT_mask = _GEN_7440 & _GEN_7189;
  assign dataArray_8_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_3_cachedata_MPORT_en = dataArray_8_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_3_cachedata_MPORT_addr = dataArray_8_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_3_cachedata_MPORT_data = dataArray_8_3[dataArray_8_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_3_MPORT_addr = replace_set;
  assign dataArray_8_3_MPORT_mask = _GEN_7440 & _GEN_7191;
  assign dataArray_8_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_4_cachedata_MPORT_en = dataArray_8_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_4_cachedata_MPORT_addr = dataArray_8_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_4_cachedata_MPORT_data = dataArray_8_4[dataArray_8_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_4_MPORT_addr = replace_set;
  assign dataArray_8_4_MPORT_mask = _GEN_7440 & _GEN_7193;
  assign dataArray_8_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_5_cachedata_MPORT_en = dataArray_8_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_5_cachedata_MPORT_addr = dataArray_8_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_5_cachedata_MPORT_data = dataArray_8_5[dataArray_8_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_5_MPORT_addr = replace_set;
  assign dataArray_8_5_MPORT_mask = _GEN_7440 & _GEN_7195;
  assign dataArray_8_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_6_cachedata_MPORT_en = dataArray_8_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_6_cachedata_MPORT_addr = dataArray_8_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_6_cachedata_MPORT_data = dataArray_8_6[dataArray_8_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_6_MPORT_addr = replace_set;
  assign dataArray_8_6_MPORT_mask = _GEN_7440 & _GEN_7197;
  assign dataArray_8_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_7_cachedata_MPORT_en = dataArray_8_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_7_cachedata_MPORT_addr = dataArray_8_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_7_cachedata_MPORT_data = dataArray_8_7[dataArray_8_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_7_MPORT_addr = replace_set;
  assign dataArray_8_7_MPORT_mask = _GEN_7440 & _GEN_7199;
  assign dataArray_8_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_8_cachedata_MPORT_en = dataArray_8_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_8_cachedata_MPORT_addr = dataArray_8_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_8_cachedata_MPORT_data = dataArray_8_8[dataArray_8_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_8_MPORT_addr = replace_set;
  assign dataArray_8_8_MPORT_mask = _GEN_7440 & _GEN_7201;
  assign dataArray_8_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_9_cachedata_MPORT_en = dataArray_8_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_9_cachedata_MPORT_addr = dataArray_8_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_9_cachedata_MPORT_data = dataArray_8_9[dataArray_8_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_9_MPORT_addr = replace_set;
  assign dataArray_8_9_MPORT_mask = _GEN_7440 & _GEN_7203;
  assign dataArray_8_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_10_cachedata_MPORT_en = dataArray_8_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_10_cachedata_MPORT_addr = dataArray_8_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_10_cachedata_MPORT_data = dataArray_8_10[dataArray_8_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_10_MPORT_addr = replace_set;
  assign dataArray_8_10_MPORT_mask = _GEN_7440 & _GEN_7205;
  assign dataArray_8_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_11_cachedata_MPORT_en = dataArray_8_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_11_cachedata_MPORT_addr = dataArray_8_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_11_cachedata_MPORT_data = dataArray_8_11[dataArray_8_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_11_MPORT_addr = replace_set;
  assign dataArray_8_11_MPORT_mask = _GEN_7440 & _GEN_7207;
  assign dataArray_8_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_12_cachedata_MPORT_en = dataArray_8_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_12_cachedata_MPORT_addr = dataArray_8_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_12_cachedata_MPORT_data = dataArray_8_12[dataArray_8_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_12_MPORT_addr = replace_set;
  assign dataArray_8_12_MPORT_mask = _GEN_7440 & _GEN_7209;
  assign dataArray_8_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_13_cachedata_MPORT_en = dataArray_8_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_13_cachedata_MPORT_addr = dataArray_8_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_13_cachedata_MPORT_data = dataArray_8_13[dataArray_8_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_13_MPORT_addr = replace_set;
  assign dataArray_8_13_MPORT_mask = _GEN_7440 & _GEN_7211;
  assign dataArray_8_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_14_cachedata_MPORT_en = dataArray_8_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_14_cachedata_MPORT_addr = dataArray_8_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_14_cachedata_MPORT_data = dataArray_8_14[dataArray_8_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_14_MPORT_addr = replace_set;
  assign dataArray_8_14_MPORT_mask = _GEN_7440 & _GEN_7213;
  assign dataArray_8_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_15_cachedata_MPORT_en = dataArray_8_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_15_cachedata_MPORT_addr = dataArray_8_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_15_cachedata_MPORT_data = dataArray_8_15[dataArray_8_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_15_MPORT_addr = replace_set;
  assign dataArray_8_15_MPORT_mask = _GEN_7440 & _GEN_7215;
  assign dataArray_8_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_0_cachedata_MPORT_en = dataArray_9_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_0_cachedata_MPORT_addr = dataArray_9_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_0_cachedata_MPORT_data = dataArray_9_0[dataArray_9_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_0_MPORT_addr = replace_set;
  assign dataArray_9_0_MPORT_mask = _GEN_7472 & _GEN_7185;
  assign dataArray_9_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_1_cachedata_MPORT_en = dataArray_9_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_1_cachedata_MPORT_addr = dataArray_9_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_1_cachedata_MPORT_data = dataArray_9_1[dataArray_9_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_1_MPORT_addr = replace_set;
  assign dataArray_9_1_MPORT_mask = _GEN_7472 & _GEN_7187;
  assign dataArray_9_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_2_cachedata_MPORT_en = dataArray_9_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_2_cachedata_MPORT_addr = dataArray_9_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_2_cachedata_MPORT_data = dataArray_9_2[dataArray_9_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_2_MPORT_addr = replace_set;
  assign dataArray_9_2_MPORT_mask = _GEN_7472 & _GEN_7189;
  assign dataArray_9_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_3_cachedata_MPORT_en = dataArray_9_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_3_cachedata_MPORT_addr = dataArray_9_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_3_cachedata_MPORT_data = dataArray_9_3[dataArray_9_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_3_MPORT_addr = replace_set;
  assign dataArray_9_3_MPORT_mask = _GEN_7472 & _GEN_7191;
  assign dataArray_9_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_4_cachedata_MPORT_en = dataArray_9_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_4_cachedata_MPORT_addr = dataArray_9_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_4_cachedata_MPORT_data = dataArray_9_4[dataArray_9_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_4_MPORT_addr = replace_set;
  assign dataArray_9_4_MPORT_mask = _GEN_7472 & _GEN_7193;
  assign dataArray_9_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_5_cachedata_MPORT_en = dataArray_9_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_5_cachedata_MPORT_addr = dataArray_9_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_5_cachedata_MPORT_data = dataArray_9_5[dataArray_9_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_5_MPORT_addr = replace_set;
  assign dataArray_9_5_MPORT_mask = _GEN_7472 & _GEN_7195;
  assign dataArray_9_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_6_cachedata_MPORT_en = dataArray_9_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_6_cachedata_MPORT_addr = dataArray_9_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_6_cachedata_MPORT_data = dataArray_9_6[dataArray_9_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_6_MPORT_addr = replace_set;
  assign dataArray_9_6_MPORT_mask = _GEN_7472 & _GEN_7197;
  assign dataArray_9_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_7_cachedata_MPORT_en = dataArray_9_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_7_cachedata_MPORT_addr = dataArray_9_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_7_cachedata_MPORT_data = dataArray_9_7[dataArray_9_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_7_MPORT_addr = replace_set;
  assign dataArray_9_7_MPORT_mask = _GEN_7472 & _GEN_7199;
  assign dataArray_9_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_8_cachedata_MPORT_en = dataArray_9_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_8_cachedata_MPORT_addr = dataArray_9_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_8_cachedata_MPORT_data = dataArray_9_8[dataArray_9_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_8_MPORT_addr = replace_set;
  assign dataArray_9_8_MPORT_mask = _GEN_7472 & _GEN_7201;
  assign dataArray_9_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_9_cachedata_MPORT_en = dataArray_9_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_9_cachedata_MPORT_addr = dataArray_9_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_9_cachedata_MPORT_data = dataArray_9_9[dataArray_9_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_9_MPORT_addr = replace_set;
  assign dataArray_9_9_MPORT_mask = _GEN_7472 & _GEN_7203;
  assign dataArray_9_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_10_cachedata_MPORT_en = dataArray_9_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_10_cachedata_MPORT_addr = dataArray_9_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_10_cachedata_MPORT_data = dataArray_9_10[dataArray_9_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_10_MPORT_addr = replace_set;
  assign dataArray_9_10_MPORT_mask = _GEN_7472 & _GEN_7205;
  assign dataArray_9_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_11_cachedata_MPORT_en = dataArray_9_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_11_cachedata_MPORT_addr = dataArray_9_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_11_cachedata_MPORT_data = dataArray_9_11[dataArray_9_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_11_MPORT_addr = replace_set;
  assign dataArray_9_11_MPORT_mask = _GEN_7472 & _GEN_7207;
  assign dataArray_9_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_12_cachedata_MPORT_en = dataArray_9_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_12_cachedata_MPORT_addr = dataArray_9_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_12_cachedata_MPORT_data = dataArray_9_12[dataArray_9_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_12_MPORT_addr = replace_set;
  assign dataArray_9_12_MPORT_mask = _GEN_7472 & _GEN_7209;
  assign dataArray_9_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_13_cachedata_MPORT_en = dataArray_9_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_13_cachedata_MPORT_addr = dataArray_9_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_13_cachedata_MPORT_data = dataArray_9_13[dataArray_9_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_13_MPORT_addr = replace_set;
  assign dataArray_9_13_MPORT_mask = _GEN_7472 & _GEN_7211;
  assign dataArray_9_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_14_cachedata_MPORT_en = dataArray_9_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_14_cachedata_MPORT_addr = dataArray_9_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_14_cachedata_MPORT_data = dataArray_9_14[dataArray_9_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_14_MPORT_addr = replace_set;
  assign dataArray_9_14_MPORT_mask = _GEN_7472 & _GEN_7213;
  assign dataArray_9_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_15_cachedata_MPORT_en = dataArray_9_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_15_cachedata_MPORT_addr = dataArray_9_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_15_cachedata_MPORT_data = dataArray_9_15[dataArray_9_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_15_MPORT_addr = replace_set;
  assign dataArray_9_15_MPORT_mask = _GEN_7472 & _GEN_7215;
  assign dataArray_9_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_0_cachedata_MPORT_en = dataArray_10_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_0_cachedata_MPORT_addr = dataArray_10_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_0_cachedata_MPORT_data = dataArray_10_0[dataArray_10_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_0_MPORT_addr = replace_set;
  assign dataArray_10_0_MPORT_mask = _GEN_7504 & _GEN_7185;
  assign dataArray_10_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_1_cachedata_MPORT_en = dataArray_10_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_1_cachedata_MPORT_addr = dataArray_10_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_1_cachedata_MPORT_data = dataArray_10_1[dataArray_10_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_1_MPORT_addr = replace_set;
  assign dataArray_10_1_MPORT_mask = _GEN_7504 & _GEN_7187;
  assign dataArray_10_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_2_cachedata_MPORT_en = dataArray_10_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_2_cachedata_MPORT_addr = dataArray_10_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_2_cachedata_MPORT_data = dataArray_10_2[dataArray_10_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_2_MPORT_addr = replace_set;
  assign dataArray_10_2_MPORT_mask = _GEN_7504 & _GEN_7189;
  assign dataArray_10_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_3_cachedata_MPORT_en = dataArray_10_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_3_cachedata_MPORT_addr = dataArray_10_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_3_cachedata_MPORT_data = dataArray_10_3[dataArray_10_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_3_MPORT_addr = replace_set;
  assign dataArray_10_3_MPORT_mask = _GEN_7504 & _GEN_7191;
  assign dataArray_10_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_4_cachedata_MPORT_en = dataArray_10_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_4_cachedata_MPORT_addr = dataArray_10_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_4_cachedata_MPORT_data = dataArray_10_4[dataArray_10_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_4_MPORT_addr = replace_set;
  assign dataArray_10_4_MPORT_mask = _GEN_7504 & _GEN_7193;
  assign dataArray_10_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_5_cachedata_MPORT_en = dataArray_10_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_5_cachedata_MPORT_addr = dataArray_10_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_5_cachedata_MPORT_data = dataArray_10_5[dataArray_10_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_5_MPORT_addr = replace_set;
  assign dataArray_10_5_MPORT_mask = _GEN_7504 & _GEN_7195;
  assign dataArray_10_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_6_cachedata_MPORT_en = dataArray_10_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_6_cachedata_MPORT_addr = dataArray_10_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_6_cachedata_MPORT_data = dataArray_10_6[dataArray_10_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_6_MPORT_addr = replace_set;
  assign dataArray_10_6_MPORT_mask = _GEN_7504 & _GEN_7197;
  assign dataArray_10_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_7_cachedata_MPORT_en = dataArray_10_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_7_cachedata_MPORT_addr = dataArray_10_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_7_cachedata_MPORT_data = dataArray_10_7[dataArray_10_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_7_MPORT_addr = replace_set;
  assign dataArray_10_7_MPORT_mask = _GEN_7504 & _GEN_7199;
  assign dataArray_10_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_8_cachedata_MPORT_en = dataArray_10_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_8_cachedata_MPORT_addr = dataArray_10_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_8_cachedata_MPORT_data = dataArray_10_8[dataArray_10_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_8_MPORT_addr = replace_set;
  assign dataArray_10_8_MPORT_mask = _GEN_7504 & _GEN_7201;
  assign dataArray_10_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_9_cachedata_MPORT_en = dataArray_10_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_9_cachedata_MPORT_addr = dataArray_10_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_9_cachedata_MPORT_data = dataArray_10_9[dataArray_10_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_9_MPORT_addr = replace_set;
  assign dataArray_10_9_MPORT_mask = _GEN_7504 & _GEN_7203;
  assign dataArray_10_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_10_cachedata_MPORT_en = dataArray_10_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_10_cachedata_MPORT_addr = dataArray_10_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_10_cachedata_MPORT_data = dataArray_10_10[dataArray_10_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_10_MPORT_addr = replace_set;
  assign dataArray_10_10_MPORT_mask = _GEN_7504 & _GEN_7205;
  assign dataArray_10_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_11_cachedata_MPORT_en = dataArray_10_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_11_cachedata_MPORT_addr = dataArray_10_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_11_cachedata_MPORT_data = dataArray_10_11[dataArray_10_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_11_MPORT_addr = replace_set;
  assign dataArray_10_11_MPORT_mask = _GEN_7504 & _GEN_7207;
  assign dataArray_10_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_12_cachedata_MPORT_en = dataArray_10_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_12_cachedata_MPORT_addr = dataArray_10_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_12_cachedata_MPORT_data = dataArray_10_12[dataArray_10_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_12_MPORT_addr = replace_set;
  assign dataArray_10_12_MPORT_mask = _GEN_7504 & _GEN_7209;
  assign dataArray_10_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_13_cachedata_MPORT_en = dataArray_10_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_13_cachedata_MPORT_addr = dataArray_10_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_13_cachedata_MPORT_data = dataArray_10_13[dataArray_10_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_13_MPORT_addr = replace_set;
  assign dataArray_10_13_MPORT_mask = _GEN_7504 & _GEN_7211;
  assign dataArray_10_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_14_cachedata_MPORT_en = dataArray_10_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_14_cachedata_MPORT_addr = dataArray_10_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_14_cachedata_MPORT_data = dataArray_10_14[dataArray_10_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_14_MPORT_addr = replace_set;
  assign dataArray_10_14_MPORT_mask = _GEN_7504 & _GEN_7213;
  assign dataArray_10_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_15_cachedata_MPORT_en = dataArray_10_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_15_cachedata_MPORT_addr = dataArray_10_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_15_cachedata_MPORT_data = dataArray_10_15[dataArray_10_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_15_MPORT_addr = replace_set;
  assign dataArray_10_15_MPORT_mask = _GEN_7504 & _GEN_7215;
  assign dataArray_10_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_0_cachedata_MPORT_en = dataArray_11_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_0_cachedata_MPORT_addr = dataArray_11_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_0_cachedata_MPORT_data = dataArray_11_0[dataArray_11_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_0_MPORT_addr = replace_set;
  assign dataArray_11_0_MPORT_mask = _GEN_7536 & _GEN_7185;
  assign dataArray_11_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_1_cachedata_MPORT_en = dataArray_11_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_1_cachedata_MPORT_addr = dataArray_11_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_1_cachedata_MPORT_data = dataArray_11_1[dataArray_11_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_1_MPORT_addr = replace_set;
  assign dataArray_11_1_MPORT_mask = _GEN_7536 & _GEN_7187;
  assign dataArray_11_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_2_cachedata_MPORT_en = dataArray_11_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_2_cachedata_MPORT_addr = dataArray_11_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_2_cachedata_MPORT_data = dataArray_11_2[dataArray_11_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_2_MPORT_addr = replace_set;
  assign dataArray_11_2_MPORT_mask = _GEN_7536 & _GEN_7189;
  assign dataArray_11_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_3_cachedata_MPORT_en = dataArray_11_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_3_cachedata_MPORT_addr = dataArray_11_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_3_cachedata_MPORT_data = dataArray_11_3[dataArray_11_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_3_MPORT_addr = replace_set;
  assign dataArray_11_3_MPORT_mask = _GEN_7536 & _GEN_7191;
  assign dataArray_11_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_4_cachedata_MPORT_en = dataArray_11_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_4_cachedata_MPORT_addr = dataArray_11_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_4_cachedata_MPORT_data = dataArray_11_4[dataArray_11_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_4_MPORT_addr = replace_set;
  assign dataArray_11_4_MPORT_mask = _GEN_7536 & _GEN_7193;
  assign dataArray_11_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_5_cachedata_MPORT_en = dataArray_11_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_5_cachedata_MPORT_addr = dataArray_11_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_5_cachedata_MPORT_data = dataArray_11_5[dataArray_11_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_5_MPORT_addr = replace_set;
  assign dataArray_11_5_MPORT_mask = _GEN_7536 & _GEN_7195;
  assign dataArray_11_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_6_cachedata_MPORT_en = dataArray_11_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_6_cachedata_MPORT_addr = dataArray_11_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_6_cachedata_MPORT_data = dataArray_11_6[dataArray_11_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_6_MPORT_addr = replace_set;
  assign dataArray_11_6_MPORT_mask = _GEN_7536 & _GEN_7197;
  assign dataArray_11_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_7_cachedata_MPORT_en = dataArray_11_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_7_cachedata_MPORT_addr = dataArray_11_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_7_cachedata_MPORT_data = dataArray_11_7[dataArray_11_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_7_MPORT_addr = replace_set;
  assign dataArray_11_7_MPORT_mask = _GEN_7536 & _GEN_7199;
  assign dataArray_11_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_8_cachedata_MPORT_en = dataArray_11_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_8_cachedata_MPORT_addr = dataArray_11_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_8_cachedata_MPORT_data = dataArray_11_8[dataArray_11_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_8_MPORT_addr = replace_set;
  assign dataArray_11_8_MPORT_mask = _GEN_7536 & _GEN_7201;
  assign dataArray_11_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_9_cachedata_MPORT_en = dataArray_11_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_9_cachedata_MPORT_addr = dataArray_11_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_9_cachedata_MPORT_data = dataArray_11_9[dataArray_11_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_9_MPORT_addr = replace_set;
  assign dataArray_11_9_MPORT_mask = _GEN_7536 & _GEN_7203;
  assign dataArray_11_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_10_cachedata_MPORT_en = dataArray_11_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_10_cachedata_MPORT_addr = dataArray_11_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_10_cachedata_MPORT_data = dataArray_11_10[dataArray_11_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_10_MPORT_addr = replace_set;
  assign dataArray_11_10_MPORT_mask = _GEN_7536 & _GEN_7205;
  assign dataArray_11_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_11_cachedata_MPORT_en = dataArray_11_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_11_cachedata_MPORT_addr = dataArray_11_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_11_cachedata_MPORT_data = dataArray_11_11[dataArray_11_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_11_MPORT_addr = replace_set;
  assign dataArray_11_11_MPORT_mask = _GEN_7536 & _GEN_7207;
  assign dataArray_11_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_12_cachedata_MPORT_en = dataArray_11_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_12_cachedata_MPORT_addr = dataArray_11_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_12_cachedata_MPORT_data = dataArray_11_12[dataArray_11_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_12_MPORT_addr = replace_set;
  assign dataArray_11_12_MPORT_mask = _GEN_7536 & _GEN_7209;
  assign dataArray_11_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_13_cachedata_MPORT_en = dataArray_11_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_13_cachedata_MPORT_addr = dataArray_11_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_13_cachedata_MPORT_data = dataArray_11_13[dataArray_11_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_13_MPORT_addr = replace_set;
  assign dataArray_11_13_MPORT_mask = _GEN_7536 & _GEN_7211;
  assign dataArray_11_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_14_cachedata_MPORT_en = dataArray_11_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_14_cachedata_MPORT_addr = dataArray_11_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_14_cachedata_MPORT_data = dataArray_11_14[dataArray_11_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_14_MPORT_addr = replace_set;
  assign dataArray_11_14_MPORT_mask = _GEN_7536 & _GEN_7213;
  assign dataArray_11_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_15_cachedata_MPORT_en = dataArray_11_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_15_cachedata_MPORT_addr = dataArray_11_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_15_cachedata_MPORT_data = dataArray_11_15[dataArray_11_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_15_MPORT_addr = replace_set;
  assign dataArray_11_15_MPORT_mask = _GEN_7536 & _GEN_7215;
  assign dataArray_11_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_0_cachedata_MPORT_en = dataArray_12_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_0_cachedata_MPORT_addr = dataArray_12_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_0_cachedata_MPORT_data = dataArray_12_0[dataArray_12_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_0_MPORT_addr = replace_set;
  assign dataArray_12_0_MPORT_mask = _GEN_7568 & _GEN_7185;
  assign dataArray_12_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_1_cachedata_MPORT_en = dataArray_12_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_1_cachedata_MPORT_addr = dataArray_12_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_1_cachedata_MPORT_data = dataArray_12_1[dataArray_12_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_1_MPORT_addr = replace_set;
  assign dataArray_12_1_MPORT_mask = _GEN_7568 & _GEN_7187;
  assign dataArray_12_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_2_cachedata_MPORT_en = dataArray_12_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_2_cachedata_MPORT_addr = dataArray_12_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_2_cachedata_MPORT_data = dataArray_12_2[dataArray_12_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_2_MPORT_addr = replace_set;
  assign dataArray_12_2_MPORT_mask = _GEN_7568 & _GEN_7189;
  assign dataArray_12_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_3_cachedata_MPORT_en = dataArray_12_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_3_cachedata_MPORT_addr = dataArray_12_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_3_cachedata_MPORT_data = dataArray_12_3[dataArray_12_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_3_MPORT_addr = replace_set;
  assign dataArray_12_3_MPORT_mask = _GEN_7568 & _GEN_7191;
  assign dataArray_12_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_4_cachedata_MPORT_en = dataArray_12_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_4_cachedata_MPORT_addr = dataArray_12_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_4_cachedata_MPORT_data = dataArray_12_4[dataArray_12_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_4_MPORT_addr = replace_set;
  assign dataArray_12_4_MPORT_mask = _GEN_7568 & _GEN_7193;
  assign dataArray_12_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_5_cachedata_MPORT_en = dataArray_12_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_5_cachedata_MPORT_addr = dataArray_12_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_5_cachedata_MPORT_data = dataArray_12_5[dataArray_12_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_5_MPORT_addr = replace_set;
  assign dataArray_12_5_MPORT_mask = _GEN_7568 & _GEN_7195;
  assign dataArray_12_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_6_cachedata_MPORT_en = dataArray_12_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_6_cachedata_MPORT_addr = dataArray_12_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_6_cachedata_MPORT_data = dataArray_12_6[dataArray_12_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_6_MPORT_addr = replace_set;
  assign dataArray_12_6_MPORT_mask = _GEN_7568 & _GEN_7197;
  assign dataArray_12_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_7_cachedata_MPORT_en = dataArray_12_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_7_cachedata_MPORT_addr = dataArray_12_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_7_cachedata_MPORT_data = dataArray_12_7[dataArray_12_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_7_MPORT_addr = replace_set;
  assign dataArray_12_7_MPORT_mask = _GEN_7568 & _GEN_7199;
  assign dataArray_12_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_8_cachedata_MPORT_en = dataArray_12_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_8_cachedata_MPORT_addr = dataArray_12_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_8_cachedata_MPORT_data = dataArray_12_8[dataArray_12_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_8_MPORT_addr = replace_set;
  assign dataArray_12_8_MPORT_mask = _GEN_7568 & _GEN_7201;
  assign dataArray_12_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_9_cachedata_MPORT_en = dataArray_12_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_9_cachedata_MPORT_addr = dataArray_12_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_9_cachedata_MPORT_data = dataArray_12_9[dataArray_12_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_9_MPORT_addr = replace_set;
  assign dataArray_12_9_MPORT_mask = _GEN_7568 & _GEN_7203;
  assign dataArray_12_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_10_cachedata_MPORT_en = dataArray_12_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_10_cachedata_MPORT_addr = dataArray_12_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_10_cachedata_MPORT_data = dataArray_12_10[dataArray_12_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_10_MPORT_addr = replace_set;
  assign dataArray_12_10_MPORT_mask = _GEN_7568 & _GEN_7205;
  assign dataArray_12_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_11_cachedata_MPORT_en = dataArray_12_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_11_cachedata_MPORT_addr = dataArray_12_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_11_cachedata_MPORT_data = dataArray_12_11[dataArray_12_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_11_MPORT_addr = replace_set;
  assign dataArray_12_11_MPORT_mask = _GEN_7568 & _GEN_7207;
  assign dataArray_12_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_12_cachedata_MPORT_en = dataArray_12_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_12_cachedata_MPORT_addr = dataArray_12_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_12_cachedata_MPORT_data = dataArray_12_12[dataArray_12_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_12_MPORT_addr = replace_set;
  assign dataArray_12_12_MPORT_mask = _GEN_7568 & _GEN_7209;
  assign dataArray_12_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_13_cachedata_MPORT_en = dataArray_12_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_13_cachedata_MPORT_addr = dataArray_12_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_13_cachedata_MPORT_data = dataArray_12_13[dataArray_12_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_13_MPORT_addr = replace_set;
  assign dataArray_12_13_MPORT_mask = _GEN_7568 & _GEN_7211;
  assign dataArray_12_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_14_cachedata_MPORT_en = dataArray_12_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_14_cachedata_MPORT_addr = dataArray_12_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_14_cachedata_MPORT_data = dataArray_12_14[dataArray_12_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_14_MPORT_addr = replace_set;
  assign dataArray_12_14_MPORT_mask = _GEN_7568 & _GEN_7213;
  assign dataArray_12_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_15_cachedata_MPORT_en = dataArray_12_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_15_cachedata_MPORT_addr = dataArray_12_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_15_cachedata_MPORT_data = dataArray_12_15[dataArray_12_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_15_MPORT_addr = replace_set;
  assign dataArray_12_15_MPORT_mask = _GEN_7568 & _GEN_7215;
  assign dataArray_12_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_0_cachedata_MPORT_en = dataArray_13_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_0_cachedata_MPORT_addr = dataArray_13_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_0_cachedata_MPORT_data = dataArray_13_0[dataArray_13_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_0_MPORT_addr = replace_set;
  assign dataArray_13_0_MPORT_mask = _GEN_7600 & _GEN_7185;
  assign dataArray_13_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_1_cachedata_MPORT_en = dataArray_13_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_1_cachedata_MPORT_addr = dataArray_13_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_1_cachedata_MPORT_data = dataArray_13_1[dataArray_13_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_1_MPORT_addr = replace_set;
  assign dataArray_13_1_MPORT_mask = _GEN_7600 & _GEN_7187;
  assign dataArray_13_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_2_cachedata_MPORT_en = dataArray_13_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_2_cachedata_MPORT_addr = dataArray_13_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_2_cachedata_MPORT_data = dataArray_13_2[dataArray_13_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_2_MPORT_addr = replace_set;
  assign dataArray_13_2_MPORT_mask = _GEN_7600 & _GEN_7189;
  assign dataArray_13_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_3_cachedata_MPORT_en = dataArray_13_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_3_cachedata_MPORT_addr = dataArray_13_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_3_cachedata_MPORT_data = dataArray_13_3[dataArray_13_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_3_MPORT_addr = replace_set;
  assign dataArray_13_3_MPORT_mask = _GEN_7600 & _GEN_7191;
  assign dataArray_13_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_4_cachedata_MPORT_en = dataArray_13_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_4_cachedata_MPORT_addr = dataArray_13_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_4_cachedata_MPORT_data = dataArray_13_4[dataArray_13_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_4_MPORT_addr = replace_set;
  assign dataArray_13_4_MPORT_mask = _GEN_7600 & _GEN_7193;
  assign dataArray_13_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_5_cachedata_MPORT_en = dataArray_13_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_5_cachedata_MPORT_addr = dataArray_13_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_5_cachedata_MPORT_data = dataArray_13_5[dataArray_13_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_5_MPORT_addr = replace_set;
  assign dataArray_13_5_MPORT_mask = _GEN_7600 & _GEN_7195;
  assign dataArray_13_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_6_cachedata_MPORT_en = dataArray_13_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_6_cachedata_MPORT_addr = dataArray_13_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_6_cachedata_MPORT_data = dataArray_13_6[dataArray_13_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_6_MPORT_addr = replace_set;
  assign dataArray_13_6_MPORT_mask = _GEN_7600 & _GEN_7197;
  assign dataArray_13_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_7_cachedata_MPORT_en = dataArray_13_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_7_cachedata_MPORT_addr = dataArray_13_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_7_cachedata_MPORT_data = dataArray_13_7[dataArray_13_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_7_MPORT_addr = replace_set;
  assign dataArray_13_7_MPORT_mask = _GEN_7600 & _GEN_7199;
  assign dataArray_13_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_8_cachedata_MPORT_en = dataArray_13_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_8_cachedata_MPORT_addr = dataArray_13_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_8_cachedata_MPORT_data = dataArray_13_8[dataArray_13_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_8_MPORT_addr = replace_set;
  assign dataArray_13_8_MPORT_mask = _GEN_7600 & _GEN_7201;
  assign dataArray_13_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_9_cachedata_MPORT_en = dataArray_13_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_9_cachedata_MPORT_addr = dataArray_13_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_9_cachedata_MPORT_data = dataArray_13_9[dataArray_13_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_9_MPORT_addr = replace_set;
  assign dataArray_13_9_MPORT_mask = _GEN_7600 & _GEN_7203;
  assign dataArray_13_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_10_cachedata_MPORT_en = dataArray_13_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_10_cachedata_MPORT_addr = dataArray_13_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_10_cachedata_MPORT_data = dataArray_13_10[dataArray_13_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_10_MPORT_addr = replace_set;
  assign dataArray_13_10_MPORT_mask = _GEN_7600 & _GEN_7205;
  assign dataArray_13_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_11_cachedata_MPORT_en = dataArray_13_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_11_cachedata_MPORT_addr = dataArray_13_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_11_cachedata_MPORT_data = dataArray_13_11[dataArray_13_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_11_MPORT_addr = replace_set;
  assign dataArray_13_11_MPORT_mask = _GEN_7600 & _GEN_7207;
  assign dataArray_13_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_12_cachedata_MPORT_en = dataArray_13_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_12_cachedata_MPORT_addr = dataArray_13_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_12_cachedata_MPORT_data = dataArray_13_12[dataArray_13_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_12_MPORT_addr = replace_set;
  assign dataArray_13_12_MPORT_mask = _GEN_7600 & _GEN_7209;
  assign dataArray_13_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_13_cachedata_MPORT_en = dataArray_13_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_13_cachedata_MPORT_addr = dataArray_13_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_13_cachedata_MPORT_data = dataArray_13_13[dataArray_13_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_13_MPORT_addr = replace_set;
  assign dataArray_13_13_MPORT_mask = _GEN_7600 & _GEN_7211;
  assign dataArray_13_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_14_cachedata_MPORT_en = dataArray_13_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_14_cachedata_MPORT_addr = dataArray_13_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_14_cachedata_MPORT_data = dataArray_13_14[dataArray_13_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_14_MPORT_addr = replace_set;
  assign dataArray_13_14_MPORT_mask = _GEN_7600 & _GEN_7213;
  assign dataArray_13_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_15_cachedata_MPORT_en = dataArray_13_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_15_cachedata_MPORT_addr = dataArray_13_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_15_cachedata_MPORT_data = dataArray_13_15[dataArray_13_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_15_MPORT_addr = replace_set;
  assign dataArray_13_15_MPORT_mask = _GEN_7600 & _GEN_7215;
  assign dataArray_13_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_0_cachedata_MPORT_en = dataArray_14_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_0_cachedata_MPORT_addr = dataArray_14_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_0_cachedata_MPORT_data = dataArray_14_0[dataArray_14_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_0_MPORT_addr = replace_set;
  assign dataArray_14_0_MPORT_mask = _GEN_7632 & _GEN_7185;
  assign dataArray_14_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_1_cachedata_MPORT_en = dataArray_14_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_1_cachedata_MPORT_addr = dataArray_14_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_1_cachedata_MPORT_data = dataArray_14_1[dataArray_14_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_1_MPORT_addr = replace_set;
  assign dataArray_14_1_MPORT_mask = _GEN_7632 & _GEN_7187;
  assign dataArray_14_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_2_cachedata_MPORT_en = dataArray_14_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_2_cachedata_MPORT_addr = dataArray_14_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_2_cachedata_MPORT_data = dataArray_14_2[dataArray_14_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_2_MPORT_addr = replace_set;
  assign dataArray_14_2_MPORT_mask = _GEN_7632 & _GEN_7189;
  assign dataArray_14_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_3_cachedata_MPORT_en = dataArray_14_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_3_cachedata_MPORT_addr = dataArray_14_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_3_cachedata_MPORT_data = dataArray_14_3[dataArray_14_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_3_MPORT_addr = replace_set;
  assign dataArray_14_3_MPORT_mask = _GEN_7632 & _GEN_7191;
  assign dataArray_14_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_4_cachedata_MPORT_en = dataArray_14_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_4_cachedata_MPORT_addr = dataArray_14_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_4_cachedata_MPORT_data = dataArray_14_4[dataArray_14_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_4_MPORT_addr = replace_set;
  assign dataArray_14_4_MPORT_mask = _GEN_7632 & _GEN_7193;
  assign dataArray_14_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_5_cachedata_MPORT_en = dataArray_14_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_5_cachedata_MPORT_addr = dataArray_14_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_5_cachedata_MPORT_data = dataArray_14_5[dataArray_14_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_5_MPORT_addr = replace_set;
  assign dataArray_14_5_MPORT_mask = _GEN_7632 & _GEN_7195;
  assign dataArray_14_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_6_cachedata_MPORT_en = dataArray_14_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_6_cachedata_MPORT_addr = dataArray_14_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_6_cachedata_MPORT_data = dataArray_14_6[dataArray_14_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_6_MPORT_addr = replace_set;
  assign dataArray_14_6_MPORT_mask = _GEN_7632 & _GEN_7197;
  assign dataArray_14_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_7_cachedata_MPORT_en = dataArray_14_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_7_cachedata_MPORT_addr = dataArray_14_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_7_cachedata_MPORT_data = dataArray_14_7[dataArray_14_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_7_MPORT_addr = replace_set;
  assign dataArray_14_7_MPORT_mask = _GEN_7632 & _GEN_7199;
  assign dataArray_14_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_8_cachedata_MPORT_en = dataArray_14_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_8_cachedata_MPORT_addr = dataArray_14_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_8_cachedata_MPORT_data = dataArray_14_8[dataArray_14_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_8_MPORT_addr = replace_set;
  assign dataArray_14_8_MPORT_mask = _GEN_7632 & _GEN_7201;
  assign dataArray_14_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_9_cachedata_MPORT_en = dataArray_14_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_9_cachedata_MPORT_addr = dataArray_14_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_9_cachedata_MPORT_data = dataArray_14_9[dataArray_14_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_9_MPORT_addr = replace_set;
  assign dataArray_14_9_MPORT_mask = _GEN_7632 & _GEN_7203;
  assign dataArray_14_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_10_cachedata_MPORT_en = dataArray_14_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_10_cachedata_MPORT_addr = dataArray_14_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_10_cachedata_MPORT_data = dataArray_14_10[dataArray_14_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_10_MPORT_addr = replace_set;
  assign dataArray_14_10_MPORT_mask = _GEN_7632 & _GEN_7205;
  assign dataArray_14_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_11_cachedata_MPORT_en = dataArray_14_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_11_cachedata_MPORT_addr = dataArray_14_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_11_cachedata_MPORT_data = dataArray_14_11[dataArray_14_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_11_MPORT_addr = replace_set;
  assign dataArray_14_11_MPORT_mask = _GEN_7632 & _GEN_7207;
  assign dataArray_14_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_12_cachedata_MPORT_en = dataArray_14_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_12_cachedata_MPORT_addr = dataArray_14_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_12_cachedata_MPORT_data = dataArray_14_12[dataArray_14_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_12_MPORT_addr = replace_set;
  assign dataArray_14_12_MPORT_mask = _GEN_7632 & _GEN_7209;
  assign dataArray_14_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_13_cachedata_MPORT_en = dataArray_14_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_13_cachedata_MPORT_addr = dataArray_14_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_13_cachedata_MPORT_data = dataArray_14_13[dataArray_14_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_13_MPORT_addr = replace_set;
  assign dataArray_14_13_MPORT_mask = _GEN_7632 & _GEN_7211;
  assign dataArray_14_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_14_cachedata_MPORT_en = dataArray_14_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_14_cachedata_MPORT_addr = dataArray_14_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_14_cachedata_MPORT_data = dataArray_14_14[dataArray_14_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_14_MPORT_addr = replace_set;
  assign dataArray_14_14_MPORT_mask = _GEN_7632 & _GEN_7213;
  assign dataArray_14_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_15_cachedata_MPORT_en = dataArray_14_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_15_cachedata_MPORT_addr = dataArray_14_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_15_cachedata_MPORT_data = dataArray_14_15[dataArray_14_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_15_MPORT_addr = replace_set;
  assign dataArray_14_15_MPORT_mask = _GEN_7632 & _GEN_7215;
  assign dataArray_14_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_0_cachedata_MPORT_en = dataArray_15_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_0_cachedata_MPORT_addr = dataArray_15_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_0_cachedata_MPORT_data = dataArray_15_0[dataArray_15_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_0_MPORT_addr = replace_set;
  assign dataArray_15_0_MPORT_mask = _GEN_7664 & _GEN_7185;
  assign dataArray_15_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_1_cachedata_MPORT_en = dataArray_15_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_1_cachedata_MPORT_addr = dataArray_15_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_1_cachedata_MPORT_data = dataArray_15_1[dataArray_15_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_1_MPORT_addr = replace_set;
  assign dataArray_15_1_MPORT_mask = _GEN_7664 & _GEN_7187;
  assign dataArray_15_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_2_cachedata_MPORT_en = dataArray_15_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_2_cachedata_MPORT_addr = dataArray_15_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_2_cachedata_MPORT_data = dataArray_15_2[dataArray_15_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_2_MPORT_addr = replace_set;
  assign dataArray_15_2_MPORT_mask = _GEN_7664 & _GEN_7189;
  assign dataArray_15_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_3_cachedata_MPORT_en = dataArray_15_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_3_cachedata_MPORT_addr = dataArray_15_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_3_cachedata_MPORT_data = dataArray_15_3[dataArray_15_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_3_MPORT_addr = replace_set;
  assign dataArray_15_3_MPORT_mask = _GEN_7664 & _GEN_7191;
  assign dataArray_15_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_4_cachedata_MPORT_en = dataArray_15_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_4_cachedata_MPORT_addr = dataArray_15_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_4_cachedata_MPORT_data = dataArray_15_4[dataArray_15_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_4_MPORT_addr = replace_set;
  assign dataArray_15_4_MPORT_mask = _GEN_7664 & _GEN_7193;
  assign dataArray_15_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_5_cachedata_MPORT_en = dataArray_15_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_5_cachedata_MPORT_addr = dataArray_15_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_5_cachedata_MPORT_data = dataArray_15_5[dataArray_15_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_5_MPORT_addr = replace_set;
  assign dataArray_15_5_MPORT_mask = _GEN_7664 & _GEN_7195;
  assign dataArray_15_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_6_cachedata_MPORT_en = dataArray_15_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_6_cachedata_MPORT_addr = dataArray_15_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_6_cachedata_MPORT_data = dataArray_15_6[dataArray_15_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_6_MPORT_addr = replace_set;
  assign dataArray_15_6_MPORT_mask = _GEN_7664 & _GEN_7197;
  assign dataArray_15_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_7_cachedata_MPORT_en = dataArray_15_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_7_cachedata_MPORT_addr = dataArray_15_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_7_cachedata_MPORT_data = dataArray_15_7[dataArray_15_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_7_MPORT_addr = replace_set;
  assign dataArray_15_7_MPORT_mask = _GEN_7664 & _GEN_7199;
  assign dataArray_15_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_8_cachedata_MPORT_en = dataArray_15_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_8_cachedata_MPORT_addr = dataArray_15_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_8_cachedata_MPORT_data = dataArray_15_8[dataArray_15_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_8_MPORT_addr = replace_set;
  assign dataArray_15_8_MPORT_mask = _GEN_7664 & _GEN_7201;
  assign dataArray_15_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_9_cachedata_MPORT_en = dataArray_15_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_9_cachedata_MPORT_addr = dataArray_15_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_9_cachedata_MPORT_data = dataArray_15_9[dataArray_15_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_9_MPORT_addr = replace_set;
  assign dataArray_15_9_MPORT_mask = _GEN_7664 & _GEN_7203;
  assign dataArray_15_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_10_cachedata_MPORT_en = dataArray_15_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_10_cachedata_MPORT_addr = dataArray_15_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_10_cachedata_MPORT_data = dataArray_15_10[dataArray_15_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_10_MPORT_addr = replace_set;
  assign dataArray_15_10_MPORT_mask = _GEN_7664 & _GEN_7205;
  assign dataArray_15_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_11_cachedata_MPORT_en = dataArray_15_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_11_cachedata_MPORT_addr = dataArray_15_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_11_cachedata_MPORT_data = dataArray_15_11[dataArray_15_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_11_MPORT_addr = replace_set;
  assign dataArray_15_11_MPORT_mask = _GEN_7664 & _GEN_7207;
  assign dataArray_15_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_12_cachedata_MPORT_en = dataArray_15_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_12_cachedata_MPORT_addr = dataArray_15_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_12_cachedata_MPORT_data = dataArray_15_12[dataArray_15_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_12_MPORT_addr = replace_set;
  assign dataArray_15_12_MPORT_mask = _GEN_7664 & _GEN_7209;
  assign dataArray_15_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_13_cachedata_MPORT_en = dataArray_15_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_13_cachedata_MPORT_addr = dataArray_15_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_13_cachedata_MPORT_data = dataArray_15_13[dataArray_15_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_13_MPORT_addr = replace_set;
  assign dataArray_15_13_MPORT_mask = _GEN_7664 & _GEN_7211;
  assign dataArray_15_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_14_cachedata_MPORT_en = dataArray_15_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_14_cachedata_MPORT_addr = dataArray_15_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_14_cachedata_MPORT_data = dataArray_15_14[dataArray_15_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_14_MPORT_addr = replace_set;
  assign dataArray_15_14_MPORT_mask = _GEN_7664 & _GEN_7213;
  assign dataArray_15_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_15_cachedata_MPORT_en = dataArray_15_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_15_cachedata_MPORT_addr = dataArray_15_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_15_cachedata_MPORT_data = dataArray_15_15[dataArray_15_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_15_MPORT_addr = replace_set;
  assign dataArray_15_15_MPORT_mask = _GEN_7664 & _GEN_7215;
  assign dataArray_15_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_0_cachedata_MPORT_en = dataArray_16_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_0_cachedata_MPORT_addr = dataArray_16_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_0_cachedata_MPORT_data = dataArray_16_0[dataArray_16_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_0_MPORT_addr = replace_set;
  assign dataArray_16_0_MPORT_mask = _GEN_7696 & _GEN_7185;
  assign dataArray_16_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_1_cachedata_MPORT_en = dataArray_16_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_1_cachedata_MPORT_addr = dataArray_16_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_1_cachedata_MPORT_data = dataArray_16_1[dataArray_16_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_1_MPORT_addr = replace_set;
  assign dataArray_16_1_MPORT_mask = _GEN_7696 & _GEN_7187;
  assign dataArray_16_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_2_cachedata_MPORT_en = dataArray_16_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_2_cachedata_MPORT_addr = dataArray_16_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_2_cachedata_MPORT_data = dataArray_16_2[dataArray_16_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_2_MPORT_addr = replace_set;
  assign dataArray_16_2_MPORT_mask = _GEN_7696 & _GEN_7189;
  assign dataArray_16_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_3_cachedata_MPORT_en = dataArray_16_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_3_cachedata_MPORT_addr = dataArray_16_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_3_cachedata_MPORT_data = dataArray_16_3[dataArray_16_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_3_MPORT_addr = replace_set;
  assign dataArray_16_3_MPORT_mask = _GEN_7696 & _GEN_7191;
  assign dataArray_16_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_4_cachedata_MPORT_en = dataArray_16_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_4_cachedata_MPORT_addr = dataArray_16_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_4_cachedata_MPORT_data = dataArray_16_4[dataArray_16_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_4_MPORT_addr = replace_set;
  assign dataArray_16_4_MPORT_mask = _GEN_7696 & _GEN_7193;
  assign dataArray_16_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_5_cachedata_MPORT_en = dataArray_16_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_5_cachedata_MPORT_addr = dataArray_16_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_5_cachedata_MPORT_data = dataArray_16_5[dataArray_16_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_5_MPORT_addr = replace_set;
  assign dataArray_16_5_MPORT_mask = _GEN_7696 & _GEN_7195;
  assign dataArray_16_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_6_cachedata_MPORT_en = dataArray_16_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_6_cachedata_MPORT_addr = dataArray_16_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_6_cachedata_MPORT_data = dataArray_16_6[dataArray_16_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_6_MPORT_addr = replace_set;
  assign dataArray_16_6_MPORT_mask = _GEN_7696 & _GEN_7197;
  assign dataArray_16_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_7_cachedata_MPORT_en = dataArray_16_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_7_cachedata_MPORT_addr = dataArray_16_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_7_cachedata_MPORT_data = dataArray_16_7[dataArray_16_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_7_MPORT_addr = replace_set;
  assign dataArray_16_7_MPORT_mask = _GEN_7696 & _GEN_7199;
  assign dataArray_16_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_8_cachedata_MPORT_en = dataArray_16_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_8_cachedata_MPORT_addr = dataArray_16_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_8_cachedata_MPORT_data = dataArray_16_8[dataArray_16_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_8_MPORT_addr = replace_set;
  assign dataArray_16_8_MPORT_mask = _GEN_7696 & _GEN_7201;
  assign dataArray_16_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_9_cachedata_MPORT_en = dataArray_16_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_9_cachedata_MPORT_addr = dataArray_16_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_9_cachedata_MPORT_data = dataArray_16_9[dataArray_16_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_9_MPORT_addr = replace_set;
  assign dataArray_16_9_MPORT_mask = _GEN_7696 & _GEN_7203;
  assign dataArray_16_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_10_cachedata_MPORT_en = dataArray_16_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_10_cachedata_MPORT_addr = dataArray_16_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_10_cachedata_MPORT_data = dataArray_16_10[dataArray_16_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_10_MPORT_addr = replace_set;
  assign dataArray_16_10_MPORT_mask = _GEN_7696 & _GEN_7205;
  assign dataArray_16_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_11_cachedata_MPORT_en = dataArray_16_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_11_cachedata_MPORT_addr = dataArray_16_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_11_cachedata_MPORT_data = dataArray_16_11[dataArray_16_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_11_MPORT_addr = replace_set;
  assign dataArray_16_11_MPORT_mask = _GEN_7696 & _GEN_7207;
  assign dataArray_16_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_12_cachedata_MPORT_en = dataArray_16_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_12_cachedata_MPORT_addr = dataArray_16_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_12_cachedata_MPORT_data = dataArray_16_12[dataArray_16_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_12_MPORT_addr = replace_set;
  assign dataArray_16_12_MPORT_mask = _GEN_7696 & _GEN_7209;
  assign dataArray_16_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_13_cachedata_MPORT_en = dataArray_16_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_13_cachedata_MPORT_addr = dataArray_16_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_13_cachedata_MPORT_data = dataArray_16_13[dataArray_16_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_13_MPORT_addr = replace_set;
  assign dataArray_16_13_MPORT_mask = _GEN_7696 & _GEN_7211;
  assign dataArray_16_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_14_cachedata_MPORT_en = dataArray_16_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_14_cachedata_MPORT_addr = dataArray_16_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_14_cachedata_MPORT_data = dataArray_16_14[dataArray_16_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_14_MPORT_addr = replace_set;
  assign dataArray_16_14_MPORT_mask = _GEN_7696 & _GEN_7213;
  assign dataArray_16_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_16_15_cachedata_MPORT_en = dataArray_16_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_16_15_cachedata_MPORT_addr = dataArray_16_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_16_15_cachedata_MPORT_data = dataArray_16_15[dataArray_16_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_16_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_16_15_MPORT_addr = replace_set;
  assign dataArray_16_15_MPORT_mask = _GEN_7696 & _GEN_7215;
  assign dataArray_16_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_0_cachedata_MPORT_en = dataArray_17_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_0_cachedata_MPORT_addr = dataArray_17_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_0_cachedata_MPORT_data = dataArray_17_0[dataArray_17_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_0_MPORT_addr = replace_set;
  assign dataArray_17_0_MPORT_mask = _GEN_7728 & _GEN_7185;
  assign dataArray_17_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_1_cachedata_MPORT_en = dataArray_17_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_1_cachedata_MPORT_addr = dataArray_17_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_1_cachedata_MPORT_data = dataArray_17_1[dataArray_17_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_1_MPORT_addr = replace_set;
  assign dataArray_17_1_MPORT_mask = _GEN_7728 & _GEN_7187;
  assign dataArray_17_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_2_cachedata_MPORT_en = dataArray_17_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_2_cachedata_MPORT_addr = dataArray_17_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_2_cachedata_MPORT_data = dataArray_17_2[dataArray_17_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_2_MPORT_addr = replace_set;
  assign dataArray_17_2_MPORT_mask = _GEN_7728 & _GEN_7189;
  assign dataArray_17_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_3_cachedata_MPORT_en = dataArray_17_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_3_cachedata_MPORT_addr = dataArray_17_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_3_cachedata_MPORT_data = dataArray_17_3[dataArray_17_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_3_MPORT_addr = replace_set;
  assign dataArray_17_3_MPORT_mask = _GEN_7728 & _GEN_7191;
  assign dataArray_17_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_4_cachedata_MPORT_en = dataArray_17_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_4_cachedata_MPORT_addr = dataArray_17_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_4_cachedata_MPORT_data = dataArray_17_4[dataArray_17_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_4_MPORT_addr = replace_set;
  assign dataArray_17_4_MPORT_mask = _GEN_7728 & _GEN_7193;
  assign dataArray_17_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_5_cachedata_MPORT_en = dataArray_17_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_5_cachedata_MPORT_addr = dataArray_17_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_5_cachedata_MPORT_data = dataArray_17_5[dataArray_17_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_5_MPORT_addr = replace_set;
  assign dataArray_17_5_MPORT_mask = _GEN_7728 & _GEN_7195;
  assign dataArray_17_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_6_cachedata_MPORT_en = dataArray_17_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_6_cachedata_MPORT_addr = dataArray_17_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_6_cachedata_MPORT_data = dataArray_17_6[dataArray_17_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_6_MPORT_addr = replace_set;
  assign dataArray_17_6_MPORT_mask = _GEN_7728 & _GEN_7197;
  assign dataArray_17_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_7_cachedata_MPORT_en = dataArray_17_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_7_cachedata_MPORT_addr = dataArray_17_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_7_cachedata_MPORT_data = dataArray_17_7[dataArray_17_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_7_MPORT_addr = replace_set;
  assign dataArray_17_7_MPORT_mask = _GEN_7728 & _GEN_7199;
  assign dataArray_17_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_8_cachedata_MPORT_en = dataArray_17_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_8_cachedata_MPORT_addr = dataArray_17_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_8_cachedata_MPORT_data = dataArray_17_8[dataArray_17_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_8_MPORT_addr = replace_set;
  assign dataArray_17_8_MPORT_mask = _GEN_7728 & _GEN_7201;
  assign dataArray_17_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_9_cachedata_MPORT_en = dataArray_17_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_9_cachedata_MPORT_addr = dataArray_17_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_9_cachedata_MPORT_data = dataArray_17_9[dataArray_17_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_9_MPORT_addr = replace_set;
  assign dataArray_17_9_MPORT_mask = _GEN_7728 & _GEN_7203;
  assign dataArray_17_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_10_cachedata_MPORT_en = dataArray_17_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_10_cachedata_MPORT_addr = dataArray_17_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_10_cachedata_MPORT_data = dataArray_17_10[dataArray_17_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_10_MPORT_addr = replace_set;
  assign dataArray_17_10_MPORT_mask = _GEN_7728 & _GEN_7205;
  assign dataArray_17_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_11_cachedata_MPORT_en = dataArray_17_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_11_cachedata_MPORT_addr = dataArray_17_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_11_cachedata_MPORT_data = dataArray_17_11[dataArray_17_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_11_MPORT_addr = replace_set;
  assign dataArray_17_11_MPORT_mask = _GEN_7728 & _GEN_7207;
  assign dataArray_17_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_12_cachedata_MPORT_en = dataArray_17_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_12_cachedata_MPORT_addr = dataArray_17_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_12_cachedata_MPORT_data = dataArray_17_12[dataArray_17_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_12_MPORT_addr = replace_set;
  assign dataArray_17_12_MPORT_mask = _GEN_7728 & _GEN_7209;
  assign dataArray_17_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_13_cachedata_MPORT_en = dataArray_17_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_13_cachedata_MPORT_addr = dataArray_17_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_13_cachedata_MPORT_data = dataArray_17_13[dataArray_17_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_13_MPORT_addr = replace_set;
  assign dataArray_17_13_MPORT_mask = _GEN_7728 & _GEN_7211;
  assign dataArray_17_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_14_cachedata_MPORT_en = dataArray_17_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_14_cachedata_MPORT_addr = dataArray_17_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_14_cachedata_MPORT_data = dataArray_17_14[dataArray_17_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_14_MPORT_addr = replace_set;
  assign dataArray_17_14_MPORT_mask = _GEN_7728 & _GEN_7213;
  assign dataArray_17_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_17_15_cachedata_MPORT_en = dataArray_17_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_17_15_cachedata_MPORT_addr = dataArray_17_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_17_15_cachedata_MPORT_data = dataArray_17_15[dataArray_17_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_17_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_17_15_MPORT_addr = replace_set;
  assign dataArray_17_15_MPORT_mask = _GEN_7728 & _GEN_7215;
  assign dataArray_17_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_0_cachedata_MPORT_en = dataArray_18_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_0_cachedata_MPORT_addr = dataArray_18_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_0_cachedata_MPORT_data = dataArray_18_0[dataArray_18_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_0_MPORT_addr = replace_set;
  assign dataArray_18_0_MPORT_mask = _GEN_7760 & _GEN_7185;
  assign dataArray_18_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_1_cachedata_MPORT_en = dataArray_18_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_1_cachedata_MPORT_addr = dataArray_18_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_1_cachedata_MPORT_data = dataArray_18_1[dataArray_18_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_1_MPORT_addr = replace_set;
  assign dataArray_18_1_MPORT_mask = _GEN_7760 & _GEN_7187;
  assign dataArray_18_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_2_cachedata_MPORT_en = dataArray_18_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_2_cachedata_MPORT_addr = dataArray_18_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_2_cachedata_MPORT_data = dataArray_18_2[dataArray_18_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_2_MPORT_addr = replace_set;
  assign dataArray_18_2_MPORT_mask = _GEN_7760 & _GEN_7189;
  assign dataArray_18_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_3_cachedata_MPORT_en = dataArray_18_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_3_cachedata_MPORT_addr = dataArray_18_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_3_cachedata_MPORT_data = dataArray_18_3[dataArray_18_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_3_MPORT_addr = replace_set;
  assign dataArray_18_3_MPORT_mask = _GEN_7760 & _GEN_7191;
  assign dataArray_18_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_4_cachedata_MPORT_en = dataArray_18_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_4_cachedata_MPORT_addr = dataArray_18_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_4_cachedata_MPORT_data = dataArray_18_4[dataArray_18_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_4_MPORT_addr = replace_set;
  assign dataArray_18_4_MPORT_mask = _GEN_7760 & _GEN_7193;
  assign dataArray_18_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_5_cachedata_MPORT_en = dataArray_18_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_5_cachedata_MPORT_addr = dataArray_18_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_5_cachedata_MPORT_data = dataArray_18_5[dataArray_18_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_5_MPORT_addr = replace_set;
  assign dataArray_18_5_MPORT_mask = _GEN_7760 & _GEN_7195;
  assign dataArray_18_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_6_cachedata_MPORT_en = dataArray_18_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_6_cachedata_MPORT_addr = dataArray_18_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_6_cachedata_MPORT_data = dataArray_18_6[dataArray_18_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_6_MPORT_addr = replace_set;
  assign dataArray_18_6_MPORT_mask = _GEN_7760 & _GEN_7197;
  assign dataArray_18_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_7_cachedata_MPORT_en = dataArray_18_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_7_cachedata_MPORT_addr = dataArray_18_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_7_cachedata_MPORT_data = dataArray_18_7[dataArray_18_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_7_MPORT_addr = replace_set;
  assign dataArray_18_7_MPORT_mask = _GEN_7760 & _GEN_7199;
  assign dataArray_18_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_8_cachedata_MPORT_en = dataArray_18_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_8_cachedata_MPORT_addr = dataArray_18_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_8_cachedata_MPORT_data = dataArray_18_8[dataArray_18_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_8_MPORT_addr = replace_set;
  assign dataArray_18_8_MPORT_mask = _GEN_7760 & _GEN_7201;
  assign dataArray_18_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_9_cachedata_MPORT_en = dataArray_18_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_9_cachedata_MPORT_addr = dataArray_18_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_9_cachedata_MPORT_data = dataArray_18_9[dataArray_18_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_9_MPORT_addr = replace_set;
  assign dataArray_18_9_MPORT_mask = _GEN_7760 & _GEN_7203;
  assign dataArray_18_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_10_cachedata_MPORT_en = dataArray_18_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_10_cachedata_MPORT_addr = dataArray_18_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_10_cachedata_MPORT_data = dataArray_18_10[dataArray_18_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_10_MPORT_addr = replace_set;
  assign dataArray_18_10_MPORT_mask = _GEN_7760 & _GEN_7205;
  assign dataArray_18_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_11_cachedata_MPORT_en = dataArray_18_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_11_cachedata_MPORT_addr = dataArray_18_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_11_cachedata_MPORT_data = dataArray_18_11[dataArray_18_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_11_MPORT_addr = replace_set;
  assign dataArray_18_11_MPORT_mask = _GEN_7760 & _GEN_7207;
  assign dataArray_18_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_12_cachedata_MPORT_en = dataArray_18_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_12_cachedata_MPORT_addr = dataArray_18_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_12_cachedata_MPORT_data = dataArray_18_12[dataArray_18_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_12_MPORT_addr = replace_set;
  assign dataArray_18_12_MPORT_mask = _GEN_7760 & _GEN_7209;
  assign dataArray_18_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_13_cachedata_MPORT_en = dataArray_18_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_13_cachedata_MPORT_addr = dataArray_18_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_13_cachedata_MPORT_data = dataArray_18_13[dataArray_18_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_13_MPORT_addr = replace_set;
  assign dataArray_18_13_MPORT_mask = _GEN_7760 & _GEN_7211;
  assign dataArray_18_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_14_cachedata_MPORT_en = dataArray_18_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_14_cachedata_MPORT_addr = dataArray_18_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_14_cachedata_MPORT_data = dataArray_18_14[dataArray_18_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_14_MPORT_addr = replace_set;
  assign dataArray_18_14_MPORT_mask = _GEN_7760 & _GEN_7213;
  assign dataArray_18_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_18_15_cachedata_MPORT_en = dataArray_18_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_18_15_cachedata_MPORT_addr = dataArray_18_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_18_15_cachedata_MPORT_data = dataArray_18_15[dataArray_18_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_18_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_18_15_MPORT_addr = replace_set;
  assign dataArray_18_15_MPORT_mask = _GEN_7760 & _GEN_7215;
  assign dataArray_18_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_0_cachedata_MPORT_en = dataArray_19_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_0_cachedata_MPORT_addr = dataArray_19_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_0_cachedata_MPORT_data = dataArray_19_0[dataArray_19_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_0_MPORT_addr = replace_set;
  assign dataArray_19_0_MPORT_mask = _GEN_7792 & _GEN_7185;
  assign dataArray_19_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_1_cachedata_MPORT_en = dataArray_19_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_1_cachedata_MPORT_addr = dataArray_19_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_1_cachedata_MPORT_data = dataArray_19_1[dataArray_19_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_1_MPORT_addr = replace_set;
  assign dataArray_19_1_MPORT_mask = _GEN_7792 & _GEN_7187;
  assign dataArray_19_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_2_cachedata_MPORT_en = dataArray_19_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_2_cachedata_MPORT_addr = dataArray_19_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_2_cachedata_MPORT_data = dataArray_19_2[dataArray_19_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_2_MPORT_addr = replace_set;
  assign dataArray_19_2_MPORT_mask = _GEN_7792 & _GEN_7189;
  assign dataArray_19_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_3_cachedata_MPORT_en = dataArray_19_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_3_cachedata_MPORT_addr = dataArray_19_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_3_cachedata_MPORT_data = dataArray_19_3[dataArray_19_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_3_MPORT_addr = replace_set;
  assign dataArray_19_3_MPORT_mask = _GEN_7792 & _GEN_7191;
  assign dataArray_19_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_4_cachedata_MPORT_en = dataArray_19_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_4_cachedata_MPORT_addr = dataArray_19_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_4_cachedata_MPORT_data = dataArray_19_4[dataArray_19_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_4_MPORT_addr = replace_set;
  assign dataArray_19_4_MPORT_mask = _GEN_7792 & _GEN_7193;
  assign dataArray_19_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_5_cachedata_MPORT_en = dataArray_19_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_5_cachedata_MPORT_addr = dataArray_19_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_5_cachedata_MPORT_data = dataArray_19_5[dataArray_19_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_5_MPORT_addr = replace_set;
  assign dataArray_19_5_MPORT_mask = _GEN_7792 & _GEN_7195;
  assign dataArray_19_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_6_cachedata_MPORT_en = dataArray_19_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_6_cachedata_MPORT_addr = dataArray_19_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_6_cachedata_MPORT_data = dataArray_19_6[dataArray_19_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_6_MPORT_addr = replace_set;
  assign dataArray_19_6_MPORT_mask = _GEN_7792 & _GEN_7197;
  assign dataArray_19_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_7_cachedata_MPORT_en = dataArray_19_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_7_cachedata_MPORT_addr = dataArray_19_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_7_cachedata_MPORT_data = dataArray_19_7[dataArray_19_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_7_MPORT_addr = replace_set;
  assign dataArray_19_7_MPORT_mask = _GEN_7792 & _GEN_7199;
  assign dataArray_19_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_8_cachedata_MPORT_en = dataArray_19_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_8_cachedata_MPORT_addr = dataArray_19_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_8_cachedata_MPORT_data = dataArray_19_8[dataArray_19_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_8_MPORT_addr = replace_set;
  assign dataArray_19_8_MPORT_mask = _GEN_7792 & _GEN_7201;
  assign dataArray_19_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_9_cachedata_MPORT_en = dataArray_19_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_9_cachedata_MPORT_addr = dataArray_19_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_9_cachedata_MPORT_data = dataArray_19_9[dataArray_19_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_9_MPORT_addr = replace_set;
  assign dataArray_19_9_MPORT_mask = _GEN_7792 & _GEN_7203;
  assign dataArray_19_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_10_cachedata_MPORT_en = dataArray_19_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_10_cachedata_MPORT_addr = dataArray_19_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_10_cachedata_MPORT_data = dataArray_19_10[dataArray_19_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_10_MPORT_addr = replace_set;
  assign dataArray_19_10_MPORT_mask = _GEN_7792 & _GEN_7205;
  assign dataArray_19_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_11_cachedata_MPORT_en = dataArray_19_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_11_cachedata_MPORT_addr = dataArray_19_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_11_cachedata_MPORT_data = dataArray_19_11[dataArray_19_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_11_MPORT_addr = replace_set;
  assign dataArray_19_11_MPORT_mask = _GEN_7792 & _GEN_7207;
  assign dataArray_19_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_12_cachedata_MPORT_en = dataArray_19_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_12_cachedata_MPORT_addr = dataArray_19_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_12_cachedata_MPORT_data = dataArray_19_12[dataArray_19_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_12_MPORT_addr = replace_set;
  assign dataArray_19_12_MPORT_mask = _GEN_7792 & _GEN_7209;
  assign dataArray_19_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_13_cachedata_MPORT_en = dataArray_19_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_13_cachedata_MPORT_addr = dataArray_19_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_13_cachedata_MPORT_data = dataArray_19_13[dataArray_19_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_13_MPORT_addr = replace_set;
  assign dataArray_19_13_MPORT_mask = _GEN_7792 & _GEN_7211;
  assign dataArray_19_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_14_cachedata_MPORT_en = dataArray_19_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_14_cachedata_MPORT_addr = dataArray_19_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_14_cachedata_MPORT_data = dataArray_19_14[dataArray_19_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_14_MPORT_addr = replace_set;
  assign dataArray_19_14_MPORT_mask = _GEN_7792 & _GEN_7213;
  assign dataArray_19_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_19_15_cachedata_MPORT_en = dataArray_19_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_19_15_cachedata_MPORT_addr = dataArray_19_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_19_15_cachedata_MPORT_data = dataArray_19_15[dataArray_19_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_19_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_19_15_MPORT_addr = replace_set;
  assign dataArray_19_15_MPORT_mask = _GEN_7792 & _GEN_7215;
  assign dataArray_19_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_0_cachedata_MPORT_en = dataArray_20_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_0_cachedata_MPORT_addr = dataArray_20_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_0_cachedata_MPORT_data = dataArray_20_0[dataArray_20_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_0_MPORT_addr = replace_set;
  assign dataArray_20_0_MPORT_mask = _GEN_7824 & _GEN_7185;
  assign dataArray_20_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_1_cachedata_MPORT_en = dataArray_20_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_1_cachedata_MPORT_addr = dataArray_20_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_1_cachedata_MPORT_data = dataArray_20_1[dataArray_20_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_1_MPORT_addr = replace_set;
  assign dataArray_20_1_MPORT_mask = _GEN_7824 & _GEN_7187;
  assign dataArray_20_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_2_cachedata_MPORT_en = dataArray_20_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_2_cachedata_MPORT_addr = dataArray_20_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_2_cachedata_MPORT_data = dataArray_20_2[dataArray_20_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_2_MPORT_addr = replace_set;
  assign dataArray_20_2_MPORT_mask = _GEN_7824 & _GEN_7189;
  assign dataArray_20_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_3_cachedata_MPORT_en = dataArray_20_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_3_cachedata_MPORT_addr = dataArray_20_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_3_cachedata_MPORT_data = dataArray_20_3[dataArray_20_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_3_MPORT_addr = replace_set;
  assign dataArray_20_3_MPORT_mask = _GEN_7824 & _GEN_7191;
  assign dataArray_20_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_4_cachedata_MPORT_en = dataArray_20_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_4_cachedata_MPORT_addr = dataArray_20_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_4_cachedata_MPORT_data = dataArray_20_4[dataArray_20_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_4_MPORT_addr = replace_set;
  assign dataArray_20_4_MPORT_mask = _GEN_7824 & _GEN_7193;
  assign dataArray_20_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_5_cachedata_MPORT_en = dataArray_20_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_5_cachedata_MPORT_addr = dataArray_20_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_5_cachedata_MPORT_data = dataArray_20_5[dataArray_20_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_5_MPORT_addr = replace_set;
  assign dataArray_20_5_MPORT_mask = _GEN_7824 & _GEN_7195;
  assign dataArray_20_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_6_cachedata_MPORT_en = dataArray_20_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_6_cachedata_MPORT_addr = dataArray_20_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_6_cachedata_MPORT_data = dataArray_20_6[dataArray_20_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_6_MPORT_addr = replace_set;
  assign dataArray_20_6_MPORT_mask = _GEN_7824 & _GEN_7197;
  assign dataArray_20_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_7_cachedata_MPORT_en = dataArray_20_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_7_cachedata_MPORT_addr = dataArray_20_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_7_cachedata_MPORT_data = dataArray_20_7[dataArray_20_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_7_MPORT_addr = replace_set;
  assign dataArray_20_7_MPORT_mask = _GEN_7824 & _GEN_7199;
  assign dataArray_20_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_8_cachedata_MPORT_en = dataArray_20_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_8_cachedata_MPORT_addr = dataArray_20_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_8_cachedata_MPORT_data = dataArray_20_8[dataArray_20_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_8_MPORT_addr = replace_set;
  assign dataArray_20_8_MPORT_mask = _GEN_7824 & _GEN_7201;
  assign dataArray_20_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_9_cachedata_MPORT_en = dataArray_20_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_9_cachedata_MPORT_addr = dataArray_20_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_9_cachedata_MPORT_data = dataArray_20_9[dataArray_20_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_9_MPORT_addr = replace_set;
  assign dataArray_20_9_MPORT_mask = _GEN_7824 & _GEN_7203;
  assign dataArray_20_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_10_cachedata_MPORT_en = dataArray_20_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_10_cachedata_MPORT_addr = dataArray_20_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_10_cachedata_MPORT_data = dataArray_20_10[dataArray_20_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_10_MPORT_addr = replace_set;
  assign dataArray_20_10_MPORT_mask = _GEN_7824 & _GEN_7205;
  assign dataArray_20_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_11_cachedata_MPORT_en = dataArray_20_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_11_cachedata_MPORT_addr = dataArray_20_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_11_cachedata_MPORT_data = dataArray_20_11[dataArray_20_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_11_MPORT_addr = replace_set;
  assign dataArray_20_11_MPORT_mask = _GEN_7824 & _GEN_7207;
  assign dataArray_20_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_12_cachedata_MPORT_en = dataArray_20_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_12_cachedata_MPORT_addr = dataArray_20_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_12_cachedata_MPORT_data = dataArray_20_12[dataArray_20_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_12_MPORT_addr = replace_set;
  assign dataArray_20_12_MPORT_mask = _GEN_7824 & _GEN_7209;
  assign dataArray_20_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_13_cachedata_MPORT_en = dataArray_20_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_13_cachedata_MPORT_addr = dataArray_20_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_13_cachedata_MPORT_data = dataArray_20_13[dataArray_20_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_13_MPORT_addr = replace_set;
  assign dataArray_20_13_MPORT_mask = _GEN_7824 & _GEN_7211;
  assign dataArray_20_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_14_cachedata_MPORT_en = dataArray_20_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_14_cachedata_MPORT_addr = dataArray_20_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_14_cachedata_MPORT_data = dataArray_20_14[dataArray_20_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_14_MPORT_addr = replace_set;
  assign dataArray_20_14_MPORT_mask = _GEN_7824 & _GEN_7213;
  assign dataArray_20_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_20_15_cachedata_MPORT_en = dataArray_20_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_20_15_cachedata_MPORT_addr = dataArray_20_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_20_15_cachedata_MPORT_data = dataArray_20_15[dataArray_20_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_20_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_20_15_MPORT_addr = replace_set;
  assign dataArray_20_15_MPORT_mask = _GEN_7824 & _GEN_7215;
  assign dataArray_20_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_0_cachedata_MPORT_en = dataArray_21_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_0_cachedata_MPORT_addr = dataArray_21_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_0_cachedata_MPORT_data = dataArray_21_0[dataArray_21_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_0_MPORT_addr = replace_set;
  assign dataArray_21_0_MPORT_mask = _GEN_7856 & _GEN_7185;
  assign dataArray_21_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_1_cachedata_MPORT_en = dataArray_21_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_1_cachedata_MPORT_addr = dataArray_21_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_1_cachedata_MPORT_data = dataArray_21_1[dataArray_21_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_1_MPORT_addr = replace_set;
  assign dataArray_21_1_MPORT_mask = _GEN_7856 & _GEN_7187;
  assign dataArray_21_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_2_cachedata_MPORT_en = dataArray_21_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_2_cachedata_MPORT_addr = dataArray_21_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_2_cachedata_MPORT_data = dataArray_21_2[dataArray_21_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_2_MPORT_addr = replace_set;
  assign dataArray_21_2_MPORT_mask = _GEN_7856 & _GEN_7189;
  assign dataArray_21_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_3_cachedata_MPORT_en = dataArray_21_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_3_cachedata_MPORT_addr = dataArray_21_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_3_cachedata_MPORT_data = dataArray_21_3[dataArray_21_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_3_MPORT_addr = replace_set;
  assign dataArray_21_3_MPORT_mask = _GEN_7856 & _GEN_7191;
  assign dataArray_21_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_4_cachedata_MPORT_en = dataArray_21_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_4_cachedata_MPORT_addr = dataArray_21_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_4_cachedata_MPORT_data = dataArray_21_4[dataArray_21_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_4_MPORT_addr = replace_set;
  assign dataArray_21_4_MPORT_mask = _GEN_7856 & _GEN_7193;
  assign dataArray_21_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_5_cachedata_MPORT_en = dataArray_21_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_5_cachedata_MPORT_addr = dataArray_21_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_5_cachedata_MPORT_data = dataArray_21_5[dataArray_21_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_5_MPORT_addr = replace_set;
  assign dataArray_21_5_MPORT_mask = _GEN_7856 & _GEN_7195;
  assign dataArray_21_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_6_cachedata_MPORT_en = dataArray_21_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_6_cachedata_MPORT_addr = dataArray_21_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_6_cachedata_MPORT_data = dataArray_21_6[dataArray_21_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_6_MPORT_addr = replace_set;
  assign dataArray_21_6_MPORT_mask = _GEN_7856 & _GEN_7197;
  assign dataArray_21_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_7_cachedata_MPORT_en = dataArray_21_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_7_cachedata_MPORT_addr = dataArray_21_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_7_cachedata_MPORT_data = dataArray_21_7[dataArray_21_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_7_MPORT_addr = replace_set;
  assign dataArray_21_7_MPORT_mask = _GEN_7856 & _GEN_7199;
  assign dataArray_21_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_8_cachedata_MPORT_en = dataArray_21_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_8_cachedata_MPORT_addr = dataArray_21_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_8_cachedata_MPORT_data = dataArray_21_8[dataArray_21_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_8_MPORT_addr = replace_set;
  assign dataArray_21_8_MPORT_mask = _GEN_7856 & _GEN_7201;
  assign dataArray_21_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_9_cachedata_MPORT_en = dataArray_21_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_9_cachedata_MPORT_addr = dataArray_21_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_9_cachedata_MPORT_data = dataArray_21_9[dataArray_21_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_9_MPORT_addr = replace_set;
  assign dataArray_21_9_MPORT_mask = _GEN_7856 & _GEN_7203;
  assign dataArray_21_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_10_cachedata_MPORT_en = dataArray_21_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_10_cachedata_MPORT_addr = dataArray_21_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_10_cachedata_MPORT_data = dataArray_21_10[dataArray_21_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_10_MPORT_addr = replace_set;
  assign dataArray_21_10_MPORT_mask = _GEN_7856 & _GEN_7205;
  assign dataArray_21_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_11_cachedata_MPORT_en = dataArray_21_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_11_cachedata_MPORT_addr = dataArray_21_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_11_cachedata_MPORT_data = dataArray_21_11[dataArray_21_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_11_MPORT_addr = replace_set;
  assign dataArray_21_11_MPORT_mask = _GEN_7856 & _GEN_7207;
  assign dataArray_21_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_12_cachedata_MPORT_en = dataArray_21_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_12_cachedata_MPORT_addr = dataArray_21_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_12_cachedata_MPORT_data = dataArray_21_12[dataArray_21_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_12_MPORT_addr = replace_set;
  assign dataArray_21_12_MPORT_mask = _GEN_7856 & _GEN_7209;
  assign dataArray_21_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_13_cachedata_MPORT_en = dataArray_21_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_13_cachedata_MPORT_addr = dataArray_21_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_13_cachedata_MPORT_data = dataArray_21_13[dataArray_21_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_13_MPORT_addr = replace_set;
  assign dataArray_21_13_MPORT_mask = _GEN_7856 & _GEN_7211;
  assign dataArray_21_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_14_cachedata_MPORT_en = dataArray_21_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_14_cachedata_MPORT_addr = dataArray_21_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_14_cachedata_MPORT_data = dataArray_21_14[dataArray_21_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_14_MPORT_addr = replace_set;
  assign dataArray_21_14_MPORT_mask = _GEN_7856 & _GEN_7213;
  assign dataArray_21_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_21_15_cachedata_MPORT_en = dataArray_21_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_21_15_cachedata_MPORT_addr = dataArray_21_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_21_15_cachedata_MPORT_data = dataArray_21_15[dataArray_21_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_21_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_21_15_MPORT_addr = replace_set;
  assign dataArray_21_15_MPORT_mask = _GEN_7856 & _GEN_7215;
  assign dataArray_21_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_0_cachedata_MPORT_en = dataArray_22_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_0_cachedata_MPORT_addr = dataArray_22_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_0_cachedata_MPORT_data = dataArray_22_0[dataArray_22_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_0_MPORT_addr = replace_set;
  assign dataArray_22_0_MPORT_mask = _GEN_7888 & _GEN_7185;
  assign dataArray_22_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_1_cachedata_MPORT_en = dataArray_22_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_1_cachedata_MPORT_addr = dataArray_22_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_1_cachedata_MPORT_data = dataArray_22_1[dataArray_22_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_1_MPORT_addr = replace_set;
  assign dataArray_22_1_MPORT_mask = _GEN_7888 & _GEN_7187;
  assign dataArray_22_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_2_cachedata_MPORT_en = dataArray_22_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_2_cachedata_MPORT_addr = dataArray_22_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_2_cachedata_MPORT_data = dataArray_22_2[dataArray_22_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_2_MPORT_addr = replace_set;
  assign dataArray_22_2_MPORT_mask = _GEN_7888 & _GEN_7189;
  assign dataArray_22_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_3_cachedata_MPORT_en = dataArray_22_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_3_cachedata_MPORT_addr = dataArray_22_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_3_cachedata_MPORT_data = dataArray_22_3[dataArray_22_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_3_MPORT_addr = replace_set;
  assign dataArray_22_3_MPORT_mask = _GEN_7888 & _GEN_7191;
  assign dataArray_22_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_4_cachedata_MPORT_en = dataArray_22_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_4_cachedata_MPORT_addr = dataArray_22_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_4_cachedata_MPORT_data = dataArray_22_4[dataArray_22_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_4_MPORT_addr = replace_set;
  assign dataArray_22_4_MPORT_mask = _GEN_7888 & _GEN_7193;
  assign dataArray_22_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_5_cachedata_MPORT_en = dataArray_22_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_5_cachedata_MPORT_addr = dataArray_22_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_5_cachedata_MPORT_data = dataArray_22_5[dataArray_22_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_5_MPORT_addr = replace_set;
  assign dataArray_22_5_MPORT_mask = _GEN_7888 & _GEN_7195;
  assign dataArray_22_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_6_cachedata_MPORT_en = dataArray_22_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_6_cachedata_MPORT_addr = dataArray_22_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_6_cachedata_MPORT_data = dataArray_22_6[dataArray_22_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_6_MPORT_addr = replace_set;
  assign dataArray_22_6_MPORT_mask = _GEN_7888 & _GEN_7197;
  assign dataArray_22_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_7_cachedata_MPORT_en = dataArray_22_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_7_cachedata_MPORT_addr = dataArray_22_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_7_cachedata_MPORT_data = dataArray_22_7[dataArray_22_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_7_MPORT_addr = replace_set;
  assign dataArray_22_7_MPORT_mask = _GEN_7888 & _GEN_7199;
  assign dataArray_22_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_8_cachedata_MPORT_en = dataArray_22_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_8_cachedata_MPORT_addr = dataArray_22_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_8_cachedata_MPORT_data = dataArray_22_8[dataArray_22_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_8_MPORT_addr = replace_set;
  assign dataArray_22_8_MPORT_mask = _GEN_7888 & _GEN_7201;
  assign dataArray_22_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_9_cachedata_MPORT_en = dataArray_22_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_9_cachedata_MPORT_addr = dataArray_22_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_9_cachedata_MPORT_data = dataArray_22_9[dataArray_22_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_9_MPORT_addr = replace_set;
  assign dataArray_22_9_MPORT_mask = _GEN_7888 & _GEN_7203;
  assign dataArray_22_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_10_cachedata_MPORT_en = dataArray_22_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_10_cachedata_MPORT_addr = dataArray_22_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_10_cachedata_MPORT_data = dataArray_22_10[dataArray_22_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_10_MPORT_addr = replace_set;
  assign dataArray_22_10_MPORT_mask = _GEN_7888 & _GEN_7205;
  assign dataArray_22_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_11_cachedata_MPORT_en = dataArray_22_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_11_cachedata_MPORT_addr = dataArray_22_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_11_cachedata_MPORT_data = dataArray_22_11[dataArray_22_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_11_MPORT_addr = replace_set;
  assign dataArray_22_11_MPORT_mask = _GEN_7888 & _GEN_7207;
  assign dataArray_22_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_12_cachedata_MPORT_en = dataArray_22_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_12_cachedata_MPORT_addr = dataArray_22_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_12_cachedata_MPORT_data = dataArray_22_12[dataArray_22_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_12_MPORT_addr = replace_set;
  assign dataArray_22_12_MPORT_mask = _GEN_7888 & _GEN_7209;
  assign dataArray_22_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_13_cachedata_MPORT_en = dataArray_22_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_13_cachedata_MPORT_addr = dataArray_22_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_13_cachedata_MPORT_data = dataArray_22_13[dataArray_22_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_13_MPORT_addr = replace_set;
  assign dataArray_22_13_MPORT_mask = _GEN_7888 & _GEN_7211;
  assign dataArray_22_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_14_cachedata_MPORT_en = dataArray_22_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_14_cachedata_MPORT_addr = dataArray_22_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_14_cachedata_MPORT_data = dataArray_22_14[dataArray_22_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_14_MPORT_addr = replace_set;
  assign dataArray_22_14_MPORT_mask = _GEN_7888 & _GEN_7213;
  assign dataArray_22_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_22_15_cachedata_MPORT_en = dataArray_22_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_22_15_cachedata_MPORT_addr = dataArray_22_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_22_15_cachedata_MPORT_data = dataArray_22_15[dataArray_22_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_22_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_22_15_MPORT_addr = replace_set;
  assign dataArray_22_15_MPORT_mask = _GEN_7888 & _GEN_7215;
  assign dataArray_22_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_0_cachedata_MPORT_en = dataArray_23_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_0_cachedata_MPORT_addr = dataArray_23_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_0_cachedata_MPORT_data = dataArray_23_0[dataArray_23_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_0_MPORT_addr = replace_set;
  assign dataArray_23_0_MPORT_mask = _GEN_7920 & _GEN_7185;
  assign dataArray_23_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_1_cachedata_MPORT_en = dataArray_23_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_1_cachedata_MPORT_addr = dataArray_23_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_1_cachedata_MPORT_data = dataArray_23_1[dataArray_23_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_1_MPORT_addr = replace_set;
  assign dataArray_23_1_MPORT_mask = _GEN_7920 & _GEN_7187;
  assign dataArray_23_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_2_cachedata_MPORT_en = dataArray_23_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_2_cachedata_MPORT_addr = dataArray_23_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_2_cachedata_MPORT_data = dataArray_23_2[dataArray_23_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_2_MPORT_addr = replace_set;
  assign dataArray_23_2_MPORT_mask = _GEN_7920 & _GEN_7189;
  assign dataArray_23_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_3_cachedata_MPORT_en = dataArray_23_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_3_cachedata_MPORT_addr = dataArray_23_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_3_cachedata_MPORT_data = dataArray_23_3[dataArray_23_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_3_MPORT_addr = replace_set;
  assign dataArray_23_3_MPORT_mask = _GEN_7920 & _GEN_7191;
  assign dataArray_23_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_4_cachedata_MPORT_en = dataArray_23_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_4_cachedata_MPORT_addr = dataArray_23_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_4_cachedata_MPORT_data = dataArray_23_4[dataArray_23_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_4_MPORT_addr = replace_set;
  assign dataArray_23_4_MPORT_mask = _GEN_7920 & _GEN_7193;
  assign dataArray_23_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_5_cachedata_MPORT_en = dataArray_23_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_5_cachedata_MPORT_addr = dataArray_23_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_5_cachedata_MPORT_data = dataArray_23_5[dataArray_23_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_5_MPORT_addr = replace_set;
  assign dataArray_23_5_MPORT_mask = _GEN_7920 & _GEN_7195;
  assign dataArray_23_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_6_cachedata_MPORT_en = dataArray_23_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_6_cachedata_MPORT_addr = dataArray_23_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_6_cachedata_MPORT_data = dataArray_23_6[dataArray_23_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_6_MPORT_addr = replace_set;
  assign dataArray_23_6_MPORT_mask = _GEN_7920 & _GEN_7197;
  assign dataArray_23_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_7_cachedata_MPORT_en = dataArray_23_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_7_cachedata_MPORT_addr = dataArray_23_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_7_cachedata_MPORT_data = dataArray_23_7[dataArray_23_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_7_MPORT_addr = replace_set;
  assign dataArray_23_7_MPORT_mask = _GEN_7920 & _GEN_7199;
  assign dataArray_23_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_8_cachedata_MPORT_en = dataArray_23_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_8_cachedata_MPORT_addr = dataArray_23_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_8_cachedata_MPORT_data = dataArray_23_8[dataArray_23_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_8_MPORT_addr = replace_set;
  assign dataArray_23_8_MPORT_mask = _GEN_7920 & _GEN_7201;
  assign dataArray_23_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_9_cachedata_MPORT_en = dataArray_23_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_9_cachedata_MPORT_addr = dataArray_23_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_9_cachedata_MPORT_data = dataArray_23_9[dataArray_23_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_9_MPORT_addr = replace_set;
  assign dataArray_23_9_MPORT_mask = _GEN_7920 & _GEN_7203;
  assign dataArray_23_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_10_cachedata_MPORT_en = dataArray_23_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_10_cachedata_MPORT_addr = dataArray_23_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_10_cachedata_MPORT_data = dataArray_23_10[dataArray_23_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_10_MPORT_addr = replace_set;
  assign dataArray_23_10_MPORT_mask = _GEN_7920 & _GEN_7205;
  assign dataArray_23_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_11_cachedata_MPORT_en = dataArray_23_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_11_cachedata_MPORT_addr = dataArray_23_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_11_cachedata_MPORT_data = dataArray_23_11[dataArray_23_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_11_MPORT_addr = replace_set;
  assign dataArray_23_11_MPORT_mask = _GEN_7920 & _GEN_7207;
  assign dataArray_23_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_12_cachedata_MPORT_en = dataArray_23_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_12_cachedata_MPORT_addr = dataArray_23_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_12_cachedata_MPORT_data = dataArray_23_12[dataArray_23_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_12_MPORT_addr = replace_set;
  assign dataArray_23_12_MPORT_mask = _GEN_7920 & _GEN_7209;
  assign dataArray_23_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_13_cachedata_MPORT_en = dataArray_23_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_13_cachedata_MPORT_addr = dataArray_23_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_13_cachedata_MPORT_data = dataArray_23_13[dataArray_23_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_13_MPORT_addr = replace_set;
  assign dataArray_23_13_MPORT_mask = _GEN_7920 & _GEN_7211;
  assign dataArray_23_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_14_cachedata_MPORT_en = dataArray_23_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_14_cachedata_MPORT_addr = dataArray_23_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_14_cachedata_MPORT_data = dataArray_23_14[dataArray_23_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_14_MPORT_addr = replace_set;
  assign dataArray_23_14_MPORT_mask = _GEN_7920 & _GEN_7213;
  assign dataArray_23_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_23_15_cachedata_MPORT_en = dataArray_23_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_23_15_cachedata_MPORT_addr = dataArray_23_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_23_15_cachedata_MPORT_data = dataArray_23_15[dataArray_23_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_23_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_23_15_MPORT_addr = replace_set;
  assign dataArray_23_15_MPORT_mask = _GEN_7920 & _GEN_7215;
  assign dataArray_23_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_0_cachedata_MPORT_en = dataArray_24_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_0_cachedata_MPORT_addr = dataArray_24_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_0_cachedata_MPORT_data = dataArray_24_0[dataArray_24_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_0_MPORT_addr = replace_set;
  assign dataArray_24_0_MPORT_mask = _GEN_7952 & _GEN_7185;
  assign dataArray_24_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_1_cachedata_MPORT_en = dataArray_24_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_1_cachedata_MPORT_addr = dataArray_24_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_1_cachedata_MPORT_data = dataArray_24_1[dataArray_24_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_1_MPORT_addr = replace_set;
  assign dataArray_24_1_MPORT_mask = _GEN_7952 & _GEN_7187;
  assign dataArray_24_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_2_cachedata_MPORT_en = dataArray_24_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_2_cachedata_MPORT_addr = dataArray_24_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_2_cachedata_MPORT_data = dataArray_24_2[dataArray_24_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_2_MPORT_addr = replace_set;
  assign dataArray_24_2_MPORT_mask = _GEN_7952 & _GEN_7189;
  assign dataArray_24_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_3_cachedata_MPORT_en = dataArray_24_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_3_cachedata_MPORT_addr = dataArray_24_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_3_cachedata_MPORT_data = dataArray_24_3[dataArray_24_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_3_MPORT_addr = replace_set;
  assign dataArray_24_3_MPORT_mask = _GEN_7952 & _GEN_7191;
  assign dataArray_24_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_4_cachedata_MPORT_en = dataArray_24_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_4_cachedata_MPORT_addr = dataArray_24_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_4_cachedata_MPORT_data = dataArray_24_4[dataArray_24_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_4_MPORT_addr = replace_set;
  assign dataArray_24_4_MPORT_mask = _GEN_7952 & _GEN_7193;
  assign dataArray_24_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_5_cachedata_MPORT_en = dataArray_24_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_5_cachedata_MPORT_addr = dataArray_24_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_5_cachedata_MPORT_data = dataArray_24_5[dataArray_24_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_5_MPORT_addr = replace_set;
  assign dataArray_24_5_MPORT_mask = _GEN_7952 & _GEN_7195;
  assign dataArray_24_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_6_cachedata_MPORT_en = dataArray_24_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_6_cachedata_MPORT_addr = dataArray_24_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_6_cachedata_MPORT_data = dataArray_24_6[dataArray_24_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_6_MPORT_addr = replace_set;
  assign dataArray_24_6_MPORT_mask = _GEN_7952 & _GEN_7197;
  assign dataArray_24_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_7_cachedata_MPORT_en = dataArray_24_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_7_cachedata_MPORT_addr = dataArray_24_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_7_cachedata_MPORT_data = dataArray_24_7[dataArray_24_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_7_MPORT_addr = replace_set;
  assign dataArray_24_7_MPORT_mask = _GEN_7952 & _GEN_7199;
  assign dataArray_24_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_8_cachedata_MPORT_en = dataArray_24_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_8_cachedata_MPORT_addr = dataArray_24_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_8_cachedata_MPORT_data = dataArray_24_8[dataArray_24_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_8_MPORT_addr = replace_set;
  assign dataArray_24_8_MPORT_mask = _GEN_7952 & _GEN_7201;
  assign dataArray_24_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_9_cachedata_MPORT_en = dataArray_24_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_9_cachedata_MPORT_addr = dataArray_24_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_9_cachedata_MPORT_data = dataArray_24_9[dataArray_24_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_9_MPORT_addr = replace_set;
  assign dataArray_24_9_MPORT_mask = _GEN_7952 & _GEN_7203;
  assign dataArray_24_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_10_cachedata_MPORT_en = dataArray_24_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_10_cachedata_MPORT_addr = dataArray_24_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_10_cachedata_MPORT_data = dataArray_24_10[dataArray_24_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_10_MPORT_addr = replace_set;
  assign dataArray_24_10_MPORT_mask = _GEN_7952 & _GEN_7205;
  assign dataArray_24_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_11_cachedata_MPORT_en = dataArray_24_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_11_cachedata_MPORT_addr = dataArray_24_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_11_cachedata_MPORT_data = dataArray_24_11[dataArray_24_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_11_MPORT_addr = replace_set;
  assign dataArray_24_11_MPORT_mask = _GEN_7952 & _GEN_7207;
  assign dataArray_24_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_12_cachedata_MPORT_en = dataArray_24_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_12_cachedata_MPORT_addr = dataArray_24_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_12_cachedata_MPORT_data = dataArray_24_12[dataArray_24_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_12_MPORT_addr = replace_set;
  assign dataArray_24_12_MPORT_mask = _GEN_7952 & _GEN_7209;
  assign dataArray_24_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_13_cachedata_MPORT_en = dataArray_24_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_13_cachedata_MPORT_addr = dataArray_24_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_13_cachedata_MPORT_data = dataArray_24_13[dataArray_24_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_13_MPORT_addr = replace_set;
  assign dataArray_24_13_MPORT_mask = _GEN_7952 & _GEN_7211;
  assign dataArray_24_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_14_cachedata_MPORT_en = dataArray_24_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_14_cachedata_MPORT_addr = dataArray_24_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_14_cachedata_MPORT_data = dataArray_24_14[dataArray_24_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_14_MPORT_addr = replace_set;
  assign dataArray_24_14_MPORT_mask = _GEN_7952 & _GEN_7213;
  assign dataArray_24_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_24_15_cachedata_MPORT_en = dataArray_24_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_24_15_cachedata_MPORT_addr = dataArray_24_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_24_15_cachedata_MPORT_data = dataArray_24_15[dataArray_24_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_24_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_24_15_MPORT_addr = replace_set;
  assign dataArray_24_15_MPORT_mask = _GEN_7952 & _GEN_7215;
  assign dataArray_24_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_0_cachedata_MPORT_en = dataArray_25_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_0_cachedata_MPORT_addr = dataArray_25_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_0_cachedata_MPORT_data = dataArray_25_0[dataArray_25_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_0_MPORT_addr = replace_set;
  assign dataArray_25_0_MPORT_mask = _GEN_7984 & _GEN_7185;
  assign dataArray_25_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_1_cachedata_MPORT_en = dataArray_25_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_1_cachedata_MPORT_addr = dataArray_25_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_1_cachedata_MPORT_data = dataArray_25_1[dataArray_25_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_1_MPORT_addr = replace_set;
  assign dataArray_25_1_MPORT_mask = _GEN_7984 & _GEN_7187;
  assign dataArray_25_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_2_cachedata_MPORT_en = dataArray_25_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_2_cachedata_MPORT_addr = dataArray_25_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_2_cachedata_MPORT_data = dataArray_25_2[dataArray_25_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_2_MPORT_addr = replace_set;
  assign dataArray_25_2_MPORT_mask = _GEN_7984 & _GEN_7189;
  assign dataArray_25_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_3_cachedata_MPORT_en = dataArray_25_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_3_cachedata_MPORT_addr = dataArray_25_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_3_cachedata_MPORT_data = dataArray_25_3[dataArray_25_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_3_MPORT_addr = replace_set;
  assign dataArray_25_3_MPORT_mask = _GEN_7984 & _GEN_7191;
  assign dataArray_25_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_4_cachedata_MPORT_en = dataArray_25_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_4_cachedata_MPORT_addr = dataArray_25_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_4_cachedata_MPORT_data = dataArray_25_4[dataArray_25_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_4_MPORT_addr = replace_set;
  assign dataArray_25_4_MPORT_mask = _GEN_7984 & _GEN_7193;
  assign dataArray_25_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_5_cachedata_MPORT_en = dataArray_25_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_5_cachedata_MPORT_addr = dataArray_25_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_5_cachedata_MPORT_data = dataArray_25_5[dataArray_25_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_5_MPORT_addr = replace_set;
  assign dataArray_25_5_MPORT_mask = _GEN_7984 & _GEN_7195;
  assign dataArray_25_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_6_cachedata_MPORT_en = dataArray_25_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_6_cachedata_MPORT_addr = dataArray_25_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_6_cachedata_MPORT_data = dataArray_25_6[dataArray_25_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_6_MPORT_addr = replace_set;
  assign dataArray_25_6_MPORT_mask = _GEN_7984 & _GEN_7197;
  assign dataArray_25_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_7_cachedata_MPORT_en = dataArray_25_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_7_cachedata_MPORT_addr = dataArray_25_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_7_cachedata_MPORT_data = dataArray_25_7[dataArray_25_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_7_MPORT_addr = replace_set;
  assign dataArray_25_7_MPORT_mask = _GEN_7984 & _GEN_7199;
  assign dataArray_25_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_8_cachedata_MPORT_en = dataArray_25_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_8_cachedata_MPORT_addr = dataArray_25_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_8_cachedata_MPORT_data = dataArray_25_8[dataArray_25_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_8_MPORT_addr = replace_set;
  assign dataArray_25_8_MPORT_mask = _GEN_7984 & _GEN_7201;
  assign dataArray_25_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_9_cachedata_MPORT_en = dataArray_25_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_9_cachedata_MPORT_addr = dataArray_25_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_9_cachedata_MPORT_data = dataArray_25_9[dataArray_25_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_9_MPORT_addr = replace_set;
  assign dataArray_25_9_MPORT_mask = _GEN_7984 & _GEN_7203;
  assign dataArray_25_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_10_cachedata_MPORT_en = dataArray_25_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_10_cachedata_MPORT_addr = dataArray_25_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_10_cachedata_MPORT_data = dataArray_25_10[dataArray_25_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_10_MPORT_addr = replace_set;
  assign dataArray_25_10_MPORT_mask = _GEN_7984 & _GEN_7205;
  assign dataArray_25_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_11_cachedata_MPORT_en = dataArray_25_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_11_cachedata_MPORT_addr = dataArray_25_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_11_cachedata_MPORT_data = dataArray_25_11[dataArray_25_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_11_MPORT_addr = replace_set;
  assign dataArray_25_11_MPORT_mask = _GEN_7984 & _GEN_7207;
  assign dataArray_25_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_12_cachedata_MPORT_en = dataArray_25_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_12_cachedata_MPORT_addr = dataArray_25_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_12_cachedata_MPORT_data = dataArray_25_12[dataArray_25_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_12_MPORT_addr = replace_set;
  assign dataArray_25_12_MPORT_mask = _GEN_7984 & _GEN_7209;
  assign dataArray_25_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_13_cachedata_MPORT_en = dataArray_25_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_13_cachedata_MPORT_addr = dataArray_25_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_13_cachedata_MPORT_data = dataArray_25_13[dataArray_25_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_13_MPORT_addr = replace_set;
  assign dataArray_25_13_MPORT_mask = _GEN_7984 & _GEN_7211;
  assign dataArray_25_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_14_cachedata_MPORT_en = dataArray_25_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_14_cachedata_MPORT_addr = dataArray_25_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_14_cachedata_MPORT_data = dataArray_25_14[dataArray_25_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_14_MPORT_addr = replace_set;
  assign dataArray_25_14_MPORT_mask = _GEN_7984 & _GEN_7213;
  assign dataArray_25_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_25_15_cachedata_MPORT_en = dataArray_25_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_25_15_cachedata_MPORT_addr = dataArray_25_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_25_15_cachedata_MPORT_data = dataArray_25_15[dataArray_25_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_25_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_25_15_MPORT_addr = replace_set;
  assign dataArray_25_15_MPORT_mask = _GEN_7984 & _GEN_7215;
  assign dataArray_25_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_0_cachedata_MPORT_en = dataArray_26_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_0_cachedata_MPORT_addr = dataArray_26_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_0_cachedata_MPORT_data = dataArray_26_0[dataArray_26_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_0_MPORT_addr = replace_set;
  assign dataArray_26_0_MPORT_mask = _GEN_8016 & _GEN_7185;
  assign dataArray_26_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_1_cachedata_MPORT_en = dataArray_26_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_1_cachedata_MPORT_addr = dataArray_26_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_1_cachedata_MPORT_data = dataArray_26_1[dataArray_26_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_1_MPORT_addr = replace_set;
  assign dataArray_26_1_MPORT_mask = _GEN_8016 & _GEN_7187;
  assign dataArray_26_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_2_cachedata_MPORT_en = dataArray_26_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_2_cachedata_MPORT_addr = dataArray_26_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_2_cachedata_MPORT_data = dataArray_26_2[dataArray_26_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_2_MPORT_addr = replace_set;
  assign dataArray_26_2_MPORT_mask = _GEN_8016 & _GEN_7189;
  assign dataArray_26_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_3_cachedata_MPORT_en = dataArray_26_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_3_cachedata_MPORT_addr = dataArray_26_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_3_cachedata_MPORT_data = dataArray_26_3[dataArray_26_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_3_MPORT_addr = replace_set;
  assign dataArray_26_3_MPORT_mask = _GEN_8016 & _GEN_7191;
  assign dataArray_26_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_4_cachedata_MPORT_en = dataArray_26_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_4_cachedata_MPORT_addr = dataArray_26_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_4_cachedata_MPORT_data = dataArray_26_4[dataArray_26_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_4_MPORT_addr = replace_set;
  assign dataArray_26_4_MPORT_mask = _GEN_8016 & _GEN_7193;
  assign dataArray_26_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_5_cachedata_MPORT_en = dataArray_26_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_5_cachedata_MPORT_addr = dataArray_26_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_5_cachedata_MPORT_data = dataArray_26_5[dataArray_26_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_5_MPORT_addr = replace_set;
  assign dataArray_26_5_MPORT_mask = _GEN_8016 & _GEN_7195;
  assign dataArray_26_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_6_cachedata_MPORT_en = dataArray_26_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_6_cachedata_MPORT_addr = dataArray_26_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_6_cachedata_MPORT_data = dataArray_26_6[dataArray_26_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_6_MPORT_addr = replace_set;
  assign dataArray_26_6_MPORT_mask = _GEN_8016 & _GEN_7197;
  assign dataArray_26_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_7_cachedata_MPORT_en = dataArray_26_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_7_cachedata_MPORT_addr = dataArray_26_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_7_cachedata_MPORT_data = dataArray_26_7[dataArray_26_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_7_MPORT_addr = replace_set;
  assign dataArray_26_7_MPORT_mask = _GEN_8016 & _GEN_7199;
  assign dataArray_26_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_8_cachedata_MPORT_en = dataArray_26_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_8_cachedata_MPORT_addr = dataArray_26_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_8_cachedata_MPORT_data = dataArray_26_8[dataArray_26_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_8_MPORT_addr = replace_set;
  assign dataArray_26_8_MPORT_mask = _GEN_8016 & _GEN_7201;
  assign dataArray_26_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_9_cachedata_MPORT_en = dataArray_26_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_9_cachedata_MPORT_addr = dataArray_26_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_9_cachedata_MPORT_data = dataArray_26_9[dataArray_26_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_9_MPORT_addr = replace_set;
  assign dataArray_26_9_MPORT_mask = _GEN_8016 & _GEN_7203;
  assign dataArray_26_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_10_cachedata_MPORT_en = dataArray_26_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_10_cachedata_MPORT_addr = dataArray_26_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_10_cachedata_MPORT_data = dataArray_26_10[dataArray_26_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_10_MPORT_addr = replace_set;
  assign dataArray_26_10_MPORT_mask = _GEN_8016 & _GEN_7205;
  assign dataArray_26_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_11_cachedata_MPORT_en = dataArray_26_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_11_cachedata_MPORT_addr = dataArray_26_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_11_cachedata_MPORT_data = dataArray_26_11[dataArray_26_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_11_MPORT_addr = replace_set;
  assign dataArray_26_11_MPORT_mask = _GEN_8016 & _GEN_7207;
  assign dataArray_26_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_12_cachedata_MPORT_en = dataArray_26_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_12_cachedata_MPORT_addr = dataArray_26_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_12_cachedata_MPORT_data = dataArray_26_12[dataArray_26_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_12_MPORT_addr = replace_set;
  assign dataArray_26_12_MPORT_mask = _GEN_8016 & _GEN_7209;
  assign dataArray_26_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_13_cachedata_MPORT_en = dataArray_26_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_13_cachedata_MPORT_addr = dataArray_26_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_13_cachedata_MPORT_data = dataArray_26_13[dataArray_26_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_13_MPORT_addr = replace_set;
  assign dataArray_26_13_MPORT_mask = _GEN_8016 & _GEN_7211;
  assign dataArray_26_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_14_cachedata_MPORT_en = dataArray_26_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_14_cachedata_MPORT_addr = dataArray_26_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_14_cachedata_MPORT_data = dataArray_26_14[dataArray_26_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_14_MPORT_addr = replace_set;
  assign dataArray_26_14_MPORT_mask = _GEN_8016 & _GEN_7213;
  assign dataArray_26_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_26_15_cachedata_MPORT_en = dataArray_26_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_26_15_cachedata_MPORT_addr = dataArray_26_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_26_15_cachedata_MPORT_data = dataArray_26_15[dataArray_26_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_26_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_26_15_MPORT_addr = replace_set;
  assign dataArray_26_15_MPORT_mask = _GEN_8016 & _GEN_7215;
  assign dataArray_26_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_0_cachedata_MPORT_en = dataArray_27_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_0_cachedata_MPORT_addr = dataArray_27_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_0_cachedata_MPORT_data = dataArray_27_0[dataArray_27_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_0_MPORT_addr = replace_set;
  assign dataArray_27_0_MPORT_mask = _GEN_8048 & _GEN_7185;
  assign dataArray_27_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_1_cachedata_MPORT_en = dataArray_27_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_1_cachedata_MPORT_addr = dataArray_27_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_1_cachedata_MPORT_data = dataArray_27_1[dataArray_27_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_1_MPORT_addr = replace_set;
  assign dataArray_27_1_MPORT_mask = _GEN_8048 & _GEN_7187;
  assign dataArray_27_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_2_cachedata_MPORT_en = dataArray_27_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_2_cachedata_MPORT_addr = dataArray_27_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_2_cachedata_MPORT_data = dataArray_27_2[dataArray_27_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_2_MPORT_addr = replace_set;
  assign dataArray_27_2_MPORT_mask = _GEN_8048 & _GEN_7189;
  assign dataArray_27_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_3_cachedata_MPORT_en = dataArray_27_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_3_cachedata_MPORT_addr = dataArray_27_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_3_cachedata_MPORT_data = dataArray_27_3[dataArray_27_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_3_MPORT_addr = replace_set;
  assign dataArray_27_3_MPORT_mask = _GEN_8048 & _GEN_7191;
  assign dataArray_27_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_4_cachedata_MPORT_en = dataArray_27_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_4_cachedata_MPORT_addr = dataArray_27_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_4_cachedata_MPORT_data = dataArray_27_4[dataArray_27_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_4_MPORT_addr = replace_set;
  assign dataArray_27_4_MPORT_mask = _GEN_8048 & _GEN_7193;
  assign dataArray_27_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_5_cachedata_MPORT_en = dataArray_27_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_5_cachedata_MPORT_addr = dataArray_27_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_5_cachedata_MPORT_data = dataArray_27_5[dataArray_27_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_5_MPORT_addr = replace_set;
  assign dataArray_27_5_MPORT_mask = _GEN_8048 & _GEN_7195;
  assign dataArray_27_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_6_cachedata_MPORT_en = dataArray_27_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_6_cachedata_MPORT_addr = dataArray_27_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_6_cachedata_MPORT_data = dataArray_27_6[dataArray_27_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_6_MPORT_addr = replace_set;
  assign dataArray_27_6_MPORT_mask = _GEN_8048 & _GEN_7197;
  assign dataArray_27_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_7_cachedata_MPORT_en = dataArray_27_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_7_cachedata_MPORT_addr = dataArray_27_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_7_cachedata_MPORT_data = dataArray_27_7[dataArray_27_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_7_MPORT_addr = replace_set;
  assign dataArray_27_7_MPORT_mask = _GEN_8048 & _GEN_7199;
  assign dataArray_27_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_8_cachedata_MPORT_en = dataArray_27_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_8_cachedata_MPORT_addr = dataArray_27_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_8_cachedata_MPORT_data = dataArray_27_8[dataArray_27_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_8_MPORT_addr = replace_set;
  assign dataArray_27_8_MPORT_mask = _GEN_8048 & _GEN_7201;
  assign dataArray_27_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_9_cachedata_MPORT_en = dataArray_27_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_9_cachedata_MPORT_addr = dataArray_27_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_9_cachedata_MPORT_data = dataArray_27_9[dataArray_27_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_9_MPORT_addr = replace_set;
  assign dataArray_27_9_MPORT_mask = _GEN_8048 & _GEN_7203;
  assign dataArray_27_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_10_cachedata_MPORT_en = dataArray_27_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_10_cachedata_MPORT_addr = dataArray_27_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_10_cachedata_MPORT_data = dataArray_27_10[dataArray_27_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_10_MPORT_addr = replace_set;
  assign dataArray_27_10_MPORT_mask = _GEN_8048 & _GEN_7205;
  assign dataArray_27_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_11_cachedata_MPORT_en = dataArray_27_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_11_cachedata_MPORT_addr = dataArray_27_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_11_cachedata_MPORT_data = dataArray_27_11[dataArray_27_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_11_MPORT_addr = replace_set;
  assign dataArray_27_11_MPORT_mask = _GEN_8048 & _GEN_7207;
  assign dataArray_27_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_12_cachedata_MPORT_en = dataArray_27_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_12_cachedata_MPORT_addr = dataArray_27_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_12_cachedata_MPORT_data = dataArray_27_12[dataArray_27_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_12_MPORT_addr = replace_set;
  assign dataArray_27_12_MPORT_mask = _GEN_8048 & _GEN_7209;
  assign dataArray_27_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_13_cachedata_MPORT_en = dataArray_27_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_13_cachedata_MPORT_addr = dataArray_27_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_13_cachedata_MPORT_data = dataArray_27_13[dataArray_27_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_13_MPORT_addr = replace_set;
  assign dataArray_27_13_MPORT_mask = _GEN_8048 & _GEN_7211;
  assign dataArray_27_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_14_cachedata_MPORT_en = dataArray_27_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_14_cachedata_MPORT_addr = dataArray_27_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_14_cachedata_MPORT_data = dataArray_27_14[dataArray_27_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_14_MPORT_addr = replace_set;
  assign dataArray_27_14_MPORT_mask = _GEN_8048 & _GEN_7213;
  assign dataArray_27_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_27_15_cachedata_MPORT_en = dataArray_27_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_27_15_cachedata_MPORT_addr = dataArray_27_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_27_15_cachedata_MPORT_data = dataArray_27_15[dataArray_27_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_27_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_27_15_MPORT_addr = replace_set;
  assign dataArray_27_15_MPORT_mask = _GEN_8048 & _GEN_7215;
  assign dataArray_27_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_0_cachedata_MPORT_en = dataArray_28_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_0_cachedata_MPORT_addr = dataArray_28_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_0_cachedata_MPORT_data = dataArray_28_0[dataArray_28_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_0_MPORT_addr = replace_set;
  assign dataArray_28_0_MPORT_mask = _GEN_8080 & _GEN_7185;
  assign dataArray_28_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_1_cachedata_MPORT_en = dataArray_28_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_1_cachedata_MPORT_addr = dataArray_28_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_1_cachedata_MPORT_data = dataArray_28_1[dataArray_28_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_1_MPORT_addr = replace_set;
  assign dataArray_28_1_MPORT_mask = _GEN_8080 & _GEN_7187;
  assign dataArray_28_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_2_cachedata_MPORT_en = dataArray_28_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_2_cachedata_MPORT_addr = dataArray_28_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_2_cachedata_MPORT_data = dataArray_28_2[dataArray_28_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_2_MPORT_addr = replace_set;
  assign dataArray_28_2_MPORT_mask = _GEN_8080 & _GEN_7189;
  assign dataArray_28_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_3_cachedata_MPORT_en = dataArray_28_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_3_cachedata_MPORT_addr = dataArray_28_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_3_cachedata_MPORT_data = dataArray_28_3[dataArray_28_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_3_MPORT_addr = replace_set;
  assign dataArray_28_3_MPORT_mask = _GEN_8080 & _GEN_7191;
  assign dataArray_28_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_4_cachedata_MPORT_en = dataArray_28_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_4_cachedata_MPORT_addr = dataArray_28_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_4_cachedata_MPORT_data = dataArray_28_4[dataArray_28_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_4_MPORT_addr = replace_set;
  assign dataArray_28_4_MPORT_mask = _GEN_8080 & _GEN_7193;
  assign dataArray_28_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_5_cachedata_MPORT_en = dataArray_28_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_5_cachedata_MPORT_addr = dataArray_28_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_5_cachedata_MPORT_data = dataArray_28_5[dataArray_28_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_5_MPORT_addr = replace_set;
  assign dataArray_28_5_MPORT_mask = _GEN_8080 & _GEN_7195;
  assign dataArray_28_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_6_cachedata_MPORT_en = dataArray_28_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_6_cachedata_MPORT_addr = dataArray_28_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_6_cachedata_MPORT_data = dataArray_28_6[dataArray_28_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_6_MPORT_addr = replace_set;
  assign dataArray_28_6_MPORT_mask = _GEN_8080 & _GEN_7197;
  assign dataArray_28_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_7_cachedata_MPORT_en = dataArray_28_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_7_cachedata_MPORT_addr = dataArray_28_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_7_cachedata_MPORT_data = dataArray_28_7[dataArray_28_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_7_MPORT_addr = replace_set;
  assign dataArray_28_7_MPORT_mask = _GEN_8080 & _GEN_7199;
  assign dataArray_28_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_8_cachedata_MPORT_en = dataArray_28_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_8_cachedata_MPORT_addr = dataArray_28_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_8_cachedata_MPORT_data = dataArray_28_8[dataArray_28_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_8_MPORT_addr = replace_set;
  assign dataArray_28_8_MPORT_mask = _GEN_8080 & _GEN_7201;
  assign dataArray_28_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_9_cachedata_MPORT_en = dataArray_28_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_9_cachedata_MPORT_addr = dataArray_28_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_9_cachedata_MPORT_data = dataArray_28_9[dataArray_28_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_9_MPORT_addr = replace_set;
  assign dataArray_28_9_MPORT_mask = _GEN_8080 & _GEN_7203;
  assign dataArray_28_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_10_cachedata_MPORT_en = dataArray_28_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_10_cachedata_MPORT_addr = dataArray_28_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_10_cachedata_MPORT_data = dataArray_28_10[dataArray_28_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_10_MPORT_addr = replace_set;
  assign dataArray_28_10_MPORT_mask = _GEN_8080 & _GEN_7205;
  assign dataArray_28_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_11_cachedata_MPORT_en = dataArray_28_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_11_cachedata_MPORT_addr = dataArray_28_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_11_cachedata_MPORT_data = dataArray_28_11[dataArray_28_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_11_MPORT_addr = replace_set;
  assign dataArray_28_11_MPORT_mask = _GEN_8080 & _GEN_7207;
  assign dataArray_28_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_12_cachedata_MPORT_en = dataArray_28_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_12_cachedata_MPORT_addr = dataArray_28_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_12_cachedata_MPORT_data = dataArray_28_12[dataArray_28_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_12_MPORT_addr = replace_set;
  assign dataArray_28_12_MPORT_mask = _GEN_8080 & _GEN_7209;
  assign dataArray_28_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_13_cachedata_MPORT_en = dataArray_28_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_13_cachedata_MPORT_addr = dataArray_28_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_13_cachedata_MPORT_data = dataArray_28_13[dataArray_28_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_13_MPORT_addr = replace_set;
  assign dataArray_28_13_MPORT_mask = _GEN_8080 & _GEN_7211;
  assign dataArray_28_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_14_cachedata_MPORT_en = dataArray_28_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_14_cachedata_MPORT_addr = dataArray_28_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_14_cachedata_MPORT_data = dataArray_28_14[dataArray_28_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_14_MPORT_addr = replace_set;
  assign dataArray_28_14_MPORT_mask = _GEN_8080 & _GEN_7213;
  assign dataArray_28_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_28_15_cachedata_MPORT_en = dataArray_28_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_28_15_cachedata_MPORT_addr = dataArray_28_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_28_15_cachedata_MPORT_data = dataArray_28_15[dataArray_28_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_28_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_28_15_MPORT_addr = replace_set;
  assign dataArray_28_15_MPORT_mask = _GEN_8080 & _GEN_7215;
  assign dataArray_28_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_0_cachedata_MPORT_en = dataArray_29_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_0_cachedata_MPORT_addr = dataArray_29_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_0_cachedata_MPORT_data = dataArray_29_0[dataArray_29_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_0_MPORT_addr = replace_set;
  assign dataArray_29_0_MPORT_mask = _GEN_8112 & _GEN_7185;
  assign dataArray_29_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_1_cachedata_MPORT_en = dataArray_29_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_1_cachedata_MPORT_addr = dataArray_29_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_1_cachedata_MPORT_data = dataArray_29_1[dataArray_29_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_1_MPORT_addr = replace_set;
  assign dataArray_29_1_MPORT_mask = _GEN_8112 & _GEN_7187;
  assign dataArray_29_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_2_cachedata_MPORT_en = dataArray_29_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_2_cachedata_MPORT_addr = dataArray_29_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_2_cachedata_MPORT_data = dataArray_29_2[dataArray_29_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_2_MPORT_addr = replace_set;
  assign dataArray_29_2_MPORT_mask = _GEN_8112 & _GEN_7189;
  assign dataArray_29_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_3_cachedata_MPORT_en = dataArray_29_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_3_cachedata_MPORT_addr = dataArray_29_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_3_cachedata_MPORT_data = dataArray_29_3[dataArray_29_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_3_MPORT_addr = replace_set;
  assign dataArray_29_3_MPORT_mask = _GEN_8112 & _GEN_7191;
  assign dataArray_29_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_4_cachedata_MPORT_en = dataArray_29_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_4_cachedata_MPORT_addr = dataArray_29_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_4_cachedata_MPORT_data = dataArray_29_4[dataArray_29_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_4_MPORT_addr = replace_set;
  assign dataArray_29_4_MPORT_mask = _GEN_8112 & _GEN_7193;
  assign dataArray_29_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_5_cachedata_MPORT_en = dataArray_29_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_5_cachedata_MPORT_addr = dataArray_29_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_5_cachedata_MPORT_data = dataArray_29_5[dataArray_29_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_5_MPORT_addr = replace_set;
  assign dataArray_29_5_MPORT_mask = _GEN_8112 & _GEN_7195;
  assign dataArray_29_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_6_cachedata_MPORT_en = dataArray_29_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_6_cachedata_MPORT_addr = dataArray_29_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_6_cachedata_MPORT_data = dataArray_29_6[dataArray_29_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_6_MPORT_addr = replace_set;
  assign dataArray_29_6_MPORT_mask = _GEN_8112 & _GEN_7197;
  assign dataArray_29_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_7_cachedata_MPORT_en = dataArray_29_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_7_cachedata_MPORT_addr = dataArray_29_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_7_cachedata_MPORT_data = dataArray_29_7[dataArray_29_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_7_MPORT_addr = replace_set;
  assign dataArray_29_7_MPORT_mask = _GEN_8112 & _GEN_7199;
  assign dataArray_29_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_8_cachedata_MPORT_en = dataArray_29_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_8_cachedata_MPORT_addr = dataArray_29_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_8_cachedata_MPORT_data = dataArray_29_8[dataArray_29_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_8_MPORT_addr = replace_set;
  assign dataArray_29_8_MPORT_mask = _GEN_8112 & _GEN_7201;
  assign dataArray_29_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_9_cachedata_MPORT_en = dataArray_29_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_9_cachedata_MPORT_addr = dataArray_29_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_9_cachedata_MPORT_data = dataArray_29_9[dataArray_29_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_9_MPORT_addr = replace_set;
  assign dataArray_29_9_MPORT_mask = _GEN_8112 & _GEN_7203;
  assign dataArray_29_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_10_cachedata_MPORT_en = dataArray_29_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_10_cachedata_MPORT_addr = dataArray_29_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_10_cachedata_MPORT_data = dataArray_29_10[dataArray_29_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_10_MPORT_addr = replace_set;
  assign dataArray_29_10_MPORT_mask = _GEN_8112 & _GEN_7205;
  assign dataArray_29_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_11_cachedata_MPORT_en = dataArray_29_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_11_cachedata_MPORT_addr = dataArray_29_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_11_cachedata_MPORT_data = dataArray_29_11[dataArray_29_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_11_MPORT_addr = replace_set;
  assign dataArray_29_11_MPORT_mask = _GEN_8112 & _GEN_7207;
  assign dataArray_29_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_12_cachedata_MPORT_en = dataArray_29_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_12_cachedata_MPORT_addr = dataArray_29_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_12_cachedata_MPORT_data = dataArray_29_12[dataArray_29_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_12_MPORT_addr = replace_set;
  assign dataArray_29_12_MPORT_mask = _GEN_8112 & _GEN_7209;
  assign dataArray_29_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_13_cachedata_MPORT_en = dataArray_29_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_13_cachedata_MPORT_addr = dataArray_29_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_13_cachedata_MPORT_data = dataArray_29_13[dataArray_29_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_13_MPORT_addr = replace_set;
  assign dataArray_29_13_MPORT_mask = _GEN_8112 & _GEN_7211;
  assign dataArray_29_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_14_cachedata_MPORT_en = dataArray_29_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_14_cachedata_MPORT_addr = dataArray_29_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_14_cachedata_MPORT_data = dataArray_29_14[dataArray_29_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_14_MPORT_addr = replace_set;
  assign dataArray_29_14_MPORT_mask = _GEN_8112 & _GEN_7213;
  assign dataArray_29_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_29_15_cachedata_MPORT_en = dataArray_29_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_29_15_cachedata_MPORT_addr = dataArray_29_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_29_15_cachedata_MPORT_data = dataArray_29_15[dataArray_29_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_29_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_29_15_MPORT_addr = replace_set;
  assign dataArray_29_15_MPORT_mask = _GEN_8112 & _GEN_7215;
  assign dataArray_29_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_0_cachedata_MPORT_en = dataArray_30_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_0_cachedata_MPORT_addr = dataArray_30_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_0_cachedata_MPORT_data = dataArray_30_0[dataArray_30_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_0_MPORT_addr = replace_set;
  assign dataArray_30_0_MPORT_mask = _GEN_8144 & _GEN_7185;
  assign dataArray_30_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_1_cachedata_MPORT_en = dataArray_30_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_1_cachedata_MPORT_addr = dataArray_30_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_1_cachedata_MPORT_data = dataArray_30_1[dataArray_30_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_1_MPORT_addr = replace_set;
  assign dataArray_30_1_MPORT_mask = _GEN_8144 & _GEN_7187;
  assign dataArray_30_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_2_cachedata_MPORT_en = dataArray_30_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_2_cachedata_MPORT_addr = dataArray_30_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_2_cachedata_MPORT_data = dataArray_30_2[dataArray_30_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_2_MPORT_addr = replace_set;
  assign dataArray_30_2_MPORT_mask = _GEN_8144 & _GEN_7189;
  assign dataArray_30_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_3_cachedata_MPORT_en = dataArray_30_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_3_cachedata_MPORT_addr = dataArray_30_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_3_cachedata_MPORT_data = dataArray_30_3[dataArray_30_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_3_MPORT_addr = replace_set;
  assign dataArray_30_3_MPORT_mask = _GEN_8144 & _GEN_7191;
  assign dataArray_30_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_4_cachedata_MPORT_en = dataArray_30_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_4_cachedata_MPORT_addr = dataArray_30_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_4_cachedata_MPORT_data = dataArray_30_4[dataArray_30_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_4_MPORT_addr = replace_set;
  assign dataArray_30_4_MPORT_mask = _GEN_8144 & _GEN_7193;
  assign dataArray_30_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_5_cachedata_MPORT_en = dataArray_30_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_5_cachedata_MPORT_addr = dataArray_30_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_5_cachedata_MPORT_data = dataArray_30_5[dataArray_30_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_5_MPORT_addr = replace_set;
  assign dataArray_30_5_MPORT_mask = _GEN_8144 & _GEN_7195;
  assign dataArray_30_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_6_cachedata_MPORT_en = dataArray_30_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_6_cachedata_MPORT_addr = dataArray_30_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_6_cachedata_MPORT_data = dataArray_30_6[dataArray_30_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_6_MPORT_addr = replace_set;
  assign dataArray_30_6_MPORT_mask = _GEN_8144 & _GEN_7197;
  assign dataArray_30_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_7_cachedata_MPORT_en = dataArray_30_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_7_cachedata_MPORT_addr = dataArray_30_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_7_cachedata_MPORT_data = dataArray_30_7[dataArray_30_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_7_MPORT_addr = replace_set;
  assign dataArray_30_7_MPORT_mask = _GEN_8144 & _GEN_7199;
  assign dataArray_30_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_8_cachedata_MPORT_en = dataArray_30_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_8_cachedata_MPORT_addr = dataArray_30_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_8_cachedata_MPORT_data = dataArray_30_8[dataArray_30_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_8_MPORT_addr = replace_set;
  assign dataArray_30_8_MPORT_mask = _GEN_8144 & _GEN_7201;
  assign dataArray_30_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_9_cachedata_MPORT_en = dataArray_30_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_9_cachedata_MPORT_addr = dataArray_30_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_9_cachedata_MPORT_data = dataArray_30_9[dataArray_30_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_9_MPORT_addr = replace_set;
  assign dataArray_30_9_MPORT_mask = _GEN_8144 & _GEN_7203;
  assign dataArray_30_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_10_cachedata_MPORT_en = dataArray_30_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_10_cachedata_MPORT_addr = dataArray_30_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_10_cachedata_MPORT_data = dataArray_30_10[dataArray_30_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_10_MPORT_addr = replace_set;
  assign dataArray_30_10_MPORT_mask = _GEN_8144 & _GEN_7205;
  assign dataArray_30_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_11_cachedata_MPORT_en = dataArray_30_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_11_cachedata_MPORT_addr = dataArray_30_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_11_cachedata_MPORT_data = dataArray_30_11[dataArray_30_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_11_MPORT_addr = replace_set;
  assign dataArray_30_11_MPORT_mask = _GEN_8144 & _GEN_7207;
  assign dataArray_30_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_12_cachedata_MPORT_en = dataArray_30_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_12_cachedata_MPORT_addr = dataArray_30_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_12_cachedata_MPORT_data = dataArray_30_12[dataArray_30_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_12_MPORT_addr = replace_set;
  assign dataArray_30_12_MPORT_mask = _GEN_8144 & _GEN_7209;
  assign dataArray_30_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_13_cachedata_MPORT_en = dataArray_30_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_13_cachedata_MPORT_addr = dataArray_30_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_13_cachedata_MPORT_data = dataArray_30_13[dataArray_30_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_13_MPORT_addr = replace_set;
  assign dataArray_30_13_MPORT_mask = _GEN_8144 & _GEN_7211;
  assign dataArray_30_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_14_cachedata_MPORT_en = dataArray_30_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_14_cachedata_MPORT_addr = dataArray_30_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_14_cachedata_MPORT_data = dataArray_30_14[dataArray_30_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_14_MPORT_addr = replace_set;
  assign dataArray_30_14_MPORT_mask = _GEN_8144 & _GEN_7213;
  assign dataArray_30_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_30_15_cachedata_MPORT_en = dataArray_30_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_30_15_cachedata_MPORT_addr = dataArray_30_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_30_15_cachedata_MPORT_data = dataArray_30_15[dataArray_30_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_30_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_30_15_MPORT_addr = replace_set;
  assign dataArray_30_15_MPORT_mask = _GEN_8144 & _GEN_7215;
  assign dataArray_30_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_0_cachedata_MPORT_en = dataArray_31_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_0_cachedata_MPORT_addr = dataArray_31_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_0_cachedata_MPORT_data = dataArray_31_0[dataArray_31_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_0_MPORT_addr = replace_set;
  assign dataArray_31_0_MPORT_mask = _GEN_8176 & _GEN_7185;
  assign dataArray_31_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_1_cachedata_MPORT_en = dataArray_31_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_1_cachedata_MPORT_addr = dataArray_31_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_1_cachedata_MPORT_data = dataArray_31_1[dataArray_31_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_1_MPORT_addr = replace_set;
  assign dataArray_31_1_MPORT_mask = _GEN_8176 & _GEN_7187;
  assign dataArray_31_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_2_cachedata_MPORT_en = dataArray_31_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_2_cachedata_MPORT_addr = dataArray_31_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_2_cachedata_MPORT_data = dataArray_31_2[dataArray_31_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_2_MPORT_addr = replace_set;
  assign dataArray_31_2_MPORT_mask = _GEN_8176 & _GEN_7189;
  assign dataArray_31_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_3_cachedata_MPORT_en = dataArray_31_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_3_cachedata_MPORT_addr = dataArray_31_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_3_cachedata_MPORT_data = dataArray_31_3[dataArray_31_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_3_MPORT_addr = replace_set;
  assign dataArray_31_3_MPORT_mask = _GEN_8176 & _GEN_7191;
  assign dataArray_31_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_4_cachedata_MPORT_en = dataArray_31_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_4_cachedata_MPORT_addr = dataArray_31_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_4_cachedata_MPORT_data = dataArray_31_4[dataArray_31_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_4_MPORT_addr = replace_set;
  assign dataArray_31_4_MPORT_mask = _GEN_8176 & _GEN_7193;
  assign dataArray_31_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_5_cachedata_MPORT_en = dataArray_31_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_5_cachedata_MPORT_addr = dataArray_31_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_5_cachedata_MPORT_data = dataArray_31_5[dataArray_31_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_5_MPORT_addr = replace_set;
  assign dataArray_31_5_MPORT_mask = _GEN_8176 & _GEN_7195;
  assign dataArray_31_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_6_cachedata_MPORT_en = dataArray_31_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_6_cachedata_MPORT_addr = dataArray_31_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_6_cachedata_MPORT_data = dataArray_31_6[dataArray_31_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_6_MPORT_addr = replace_set;
  assign dataArray_31_6_MPORT_mask = _GEN_8176 & _GEN_7197;
  assign dataArray_31_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_7_cachedata_MPORT_en = dataArray_31_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_7_cachedata_MPORT_addr = dataArray_31_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_7_cachedata_MPORT_data = dataArray_31_7[dataArray_31_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_7_MPORT_addr = replace_set;
  assign dataArray_31_7_MPORT_mask = _GEN_8176 & _GEN_7199;
  assign dataArray_31_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_8_cachedata_MPORT_en = dataArray_31_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_8_cachedata_MPORT_addr = dataArray_31_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_8_cachedata_MPORT_data = dataArray_31_8[dataArray_31_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_8_MPORT_addr = replace_set;
  assign dataArray_31_8_MPORT_mask = _GEN_8176 & _GEN_7201;
  assign dataArray_31_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_9_cachedata_MPORT_en = dataArray_31_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_9_cachedata_MPORT_addr = dataArray_31_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_9_cachedata_MPORT_data = dataArray_31_9[dataArray_31_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_9_MPORT_addr = replace_set;
  assign dataArray_31_9_MPORT_mask = _GEN_8176 & _GEN_7203;
  assign dataArray_31_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_10_cachedata_MPORT_en = dataArray_31_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_10_cachedata_MPORT_addr = dataArray_31_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_10_cachedata_MPORT_data = dataArray_31_10[dataArray_31_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_10_MPORT_addr = replace_set;
  assign dataArray_31_10_MPORT_mask = _GEN_8176 & _GEN_7205;
  assign dataArray_31_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_11_cachedata_MPORT_en = dataArray_31_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_11_cachedata_MPORT_addr = dataArray_31_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_11_cachedata_MPORT_data = dataArray_31_11[dataArray_31_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_11_MPORT_addr = replace_set;
  assign dataArray_31_11_MPORT_mask = _GEN_8176 & _GEN_7207;
  assign dataArray_31_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_12_cachedata_MPORT_en = dataArray_31_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_12_cachedata_MPORT_addr = dataArray_31_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_12_cachedata_MPORT_data = dataArray_31_12[dataArray_31_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_12_MPORT_addr = replace_set;
  assign dataArray_31_12_MPORT_mask = _GEN_8176 & _GEN_7209;
  assign dataArray_31_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_13_cachedata_MPORT_en = dataArray_31_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_13_cachedata_MPORT_addr = dataArray_31_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_13_cachedata_MPORT_data = dataArray_31_13[dataArray_31_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_13_MPORT_addr = replace_set;
  assign dataArray_31_13_MPORT_mask = _GEN_8176 & _GEN_7211;
  assign dataArray_31_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_14_cachedata_MPORT_en = dataArray_31_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_14_cachedata_MPORT_addr = dataArray_31_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_14_cachedata_MPORT_data = dataArray_31_14[dataArray_31_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_14_MPORT_addr = replace_set;
  assign dataArray_31_14_MPORT_mask = _GEN_8176 & _GEN_7213;
  assign dataArray_31_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_31_15_cachedata_MPORT_en = dataArray_31_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_31_15_cachedata_MPORT_addr = dataArray_31_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_31_15_cachedata_MPORT_data = dataArray_31_15[dataArray_31_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_31_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_31_15_MPORT_addr = replace_set;
  assign dataArray_31_15_MPORT_mask = _GEN_8176 & _GEN_7215;
  assign dataArray_31_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_0_cachedata_MPORT_en = dataArray_32_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_0_cachedata_MPORT_addr = dataArray_32_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_0_cachedata_MPORT_data = dataArray_32_0[dataArray_32_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_0_MPORT_addr = replace_set;
  assign dataArray_32_0_MPORT_mask = _GEN_8208 & _GEN_7185;
  assign dataArray_32_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_1_cachedata_MPORT_en = dataArray_32_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_1_cachedata_MPORT_addr = dataArray_32_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_1_cachedata_MPORT_data = dataArray_32_1[dataArray_32_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_1_MPORT_addr = replace_set;
  assign dataArray_32_1_MPORT_mask = _GEN_8208 & _GEN_7187;
  assign dataArray_32_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_2_cachedata_MPORT_en = dataArray_32_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_2_cachedata_MPORT_addr = dataArray_32_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_2_cachedata_MPORT_data = dataArray_32_2[dataArray_32_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_2_MPORT_addr = replace_set;
  assign dataArray_32_2_MPORT_mask = _GEN_8208 & _GEN_7189;
  assign dataArray_32_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_3_cachedata_MPORT_en = dataArray_32_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_3_cachedata_MPORT_addr = dataArray_32_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_3_cachedata_MPORT_data = dataArray_32_3[dataArray_32_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_3_MPORT_addr = replace_set;
  assign dataArray_32_3_MPORT_mask = _GEN_8208 & _GEN_7191;
  assign dataArray_32_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_4_cachedata_MPORT_en = dataArray_32_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_4_cachedata_MPORT_addr = dataArray_32_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_4_cachedata_MPORT_data = dataArray_32_4[dataArray_32_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_4_MPORT_addr = replace_set;
  assign dataArray_32_4_MPORT_mask = _GEN_8208 & _GEN_7193;
  assign dataArray_32_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_5_cachedata_MPORT_en = dataArray_32_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_5_cachedata_MPORT_addr = dataArray_32_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_5_cachedata_MPORT_data = dataArray_32_5[dataArray_32_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_5_MPORT_addr = replace_set;
  assign dataArray_32_5_MPORT_mask = _GEN_8208 & _GEN_7195;
  assign dataArray_32_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_6_cachedata_MPORT_en = dataArray_32_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_6_cachedata_MPORT_addr = dataArray_32_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_6_cachedata_MPORT_data = dataArray_32_6[dataArray_32_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_6_MPORT_addr = replace_set;
  assign dataArray_32_6_MPORT_mask = _GEN_8208 & _GEN_7197;
  assign dataArray_32_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_7_cachedata_MPORT_en = dataArray_32_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_7_cachedata_MPORT_addr = dataArray_32_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_7_cachedata_MPORT_data = dataArray_32_7[dataArray_32_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_7_MPORT_addr = replace_set;
  assign dataArray_32_7_MPORT_mask = _GEN_8208 & _GEN_7199;
  assign dataArray_32_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_8_cachedata_MPORT_en = dataArray_32_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_8_cachedata_MPORT_addr = dataArray_32_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_8_cachedata_MPORT_data = dataArray_32_8[dataArray_32_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_8_MPORT_addr = replace_set;
  assign dataArray_32_8_MPORT_mask = _GEN_8208 & _GEN_7201;
  assign dataArray_32_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_9_cachedata_MPORT_en = dataArray_32_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_9_cachedata_MPORT_addr = dataArray_32_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_9_cachedata_MPORT_data = dataArray_32_9[dataArray_32_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_9_MPORT_addr = replace_set;
  assign dataArray_32_9_MPORT_mask = _GEN_8208 & _GEN_7203;
  assign dataArray_32_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_10_cachedata_MPORT_en = dataArray_32_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_10_cachedata_MPORT_addr = dataArray_32_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_10_cachedata_MPORT_data = dataArray_32_10[dataArray_32_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_10_MPORT_addr = replace_set;
  assign dataArray_32_10_MPORT_mask = _GEN_8208 & _GEN_7205;
  assign dataArray_32_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_11_cachedata_MPORT_en = dataArray_32_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_11_cachedata_MPORT_addr = dataArray_32_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_11_cachedata_MPORT_data = dataArray_32_11[dataArray_32_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_11_MPORT_addr = replace_set;
  assign dataArray_32_11_MPORT_mask = _GEN_8208 & _GEN_7207;
  assign dataArray_32_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_12_cachedata_MPORT_en = dataArray_32_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_12_cachedata_MPORT_addr = dataArray_32_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_12_cachedata_MPORT_data = dataArray_32_12[dataArray_32_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_12_MPORT_addr = replace_set;
  assign dataArray_32_12_MPORT_mask = _GEN_8208 & _GEN_7209;
  assign dataArray_32_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_13_cachedata_MPORT_en = dataArray_32_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_13_cachedata_MPORT_addr = dataArray_32_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_13_cachedata_MPORT_data = dataArray_32_13[dataArray_32_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_13_MPORT_addr = replace_set;
  assign dataArray_32_13_MPORT_mask = _GEN_8208 & _GEN_7211;
  assign dataArray_32_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_14_cachedata_MPORT_en = dataArray_32_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_14_cachedata_MPORT_addr = dataArray_32_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_14_cachedata_MPORT_data = dataArray_32_14[dataArray_32_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_14_MPORT_addr = replace_set;
  assign dataArray_32_14_MPORT_mask = _GEN_8208 & _GEN_7213;
  assign dataArray_32_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_32_15_cachedata_MPORT_en = dataArray_32_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_32_15_cachedata_MPORT_addr = dataArray_32_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_32_15_cachedata_MPORT_data = dataArray_32_15[dataArray_32_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_32_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_32_15_MPORT_addr = replace_set;
  assign dataArray_32_15_MPORT_mask = _GEN_8208 & _GEN_7215;
  assign dataArray_32_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_0_cachedata_MPORT_en = dataArray_33_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_0_cachedata_MPORT_addr = dataArray_33_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_0_cachedata_MPORT_data = dataArray_33_0[dataArray_33_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_0_MPORT_addr = replace_set;
  assign dataArray_33_0_MPORT_mask = _GEN_8240 & _GEN_7185;
  assign dataArray_33_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_1_cachedata_MPORT_en = dataArray_33_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_1_cachedata_MPORT_addr = dataArray_33_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_1_cachedata_MPORT_data = dataArray_33_1[dataArray_33_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_1_MPORT_addr = replace_set;
  assign dataArray_33_1_MPORT_mask = _GEN_8240 & _GEN_7187;
  assign dataArray_33_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_2_cachedata_MPORT_en = dataArray_33_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_2_cachedata_MPORT_addr = dataArray_33_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_2_cachedata_MPORT_data = dataArray_33_2[dataArray_33_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_2_MPORT_addr = replace_set;
  assign dataArray_33_2_MPORT_mask = _GEN_8240 & _GEN_7189;
  assign dataArray_33_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_3_cachedata_MPORT_en = dataArray_33_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_3_cachedata_MPORT_addr = dataArray_33_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_3_cachedata_MPORT_data = dataArray_33_3[dataArray_33_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_3_MPORT_addr = replace_set;
  assign dataArray_33_3_MPORT_mask = _GEN_8240 & _GEN_7191;
  assign dataArray_33_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_4_cachedata_MPORT_en = dataArray_33_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_4_cachedata_MPORT_addr = dataArray_33_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_4_cachedata_MPORT_data = dataArray_33_4[dataArray_33_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_4_MPORT_addr = replace_set;
  assign dataArray_33_4_MPORT_mask = _GEN_8240 & _GEN_7193;
  assign dataArray_33_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_5_cachedata_MPORT_en = dataArray_33_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_5_cachedata_MPORT_addr = dataArray_33_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_5_cachedata_MPORT_data = dataArray_33_5[dataArray_33_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_5_MPORT_addr = replace_set;
  assign dataArray_33_5_MPORT_mask = _GEN_8240 & _GEN_7195;
  assign dataArray_33_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_6_cachedata_MPORT_en = dataArray_33_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_6_cachedata_MPORT_addr = dataArray_33_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_6_cachedata_MPORT_data = dataArray_33_6[dataArray_33_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_6_MPORT_addr = replace_set;
  assign dataArray_33_6_MPORT_mask = _GEN_8240 & _GEN_7197;
  assign dataArray_33_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_7_cachedata_MPORT_en = dataArray_33_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_7_cachedata_MPORT_addr = dataArray_33_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_7_cachedata_MPORT_data = dataArray_33_7[dataArray_33_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_7_MPORT_addr = replace_set;
  assign dataArray_33_7_MPORT_mask = _GEN_8240 & _GEN_7199;
  assign dataArray_33_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_8_cachedata_MPORT_en = dataArray_33_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_8_cachedata_MPORT_addr = dataArray_33_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_8_cachedata_MPORT_data = dataArray_33_8[dataArray_33_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_8_MPORT_addr = replace_set;
  assign dataArray_33_8_MPORT_mask = _GEN_8240 & _GEN_7201;
  assign dataArray_33_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_9_cachedata_MPORT_en = dataArray_33_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_9_cachedata_MPORT_addr = dataArray_33_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_9_cachedata_MPORT_data = dataArray_33_9[dataArray_33_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_9_MPORT_addr = replace_set;
  assign dataArray_33_9_MPORT_mask = _GEN_8240 & _GEN_7203;
  assign dataArray_33_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_10_cachedata_MPORT_en = dataArray_33_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_10_cachedata_MPORT_addr = dataArray_33_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_10_cachedata_MPORT_data = dataArray_33_10[dataArray_33_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_10_MPORT_addr = replace_set;
  assign dataArray_33_10_MPORT_mask = _GEN_8240 & _GEN_7205;
  assign dataArray_33_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_11_cachedata_MPORT_en = dataArray_33_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_11_cachedata_MPORT_addr = dataArray_33_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_11_cachedata_MPORT_data = dataArray_33_11[dataArray_33_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_11_MPORT_addr = replace_set;
  assign dataArray_33_11_MPORT_mask = _GEN_8240 & _GEN_7207;
  assign dataArray_33_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_12_cachedata_MPORT_en = dataArray_33_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_12_cachedata_MPORT_addr = dataArray_33_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_12_cachedata_MPORT_data = dataArray_33_12[dataArray_33_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_12_MPORT_addr = replace_set;
  assign dataArray_33_12_MPORT_mask = _GEN_8240 & _GEN_7209;
  assign dataArray_33_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_13_cachedata_MPORT_en = dataArray_33_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_13_cachedata_MPORT_addr = dataArray_33_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_13_cachedata_MPORT_data = dataArray_33_13[dataArray_33_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_13_MPORT_addr = replace_set;
  assign dataArray_33_13_MPORT_mask = _GEN_8240 & _GEN_7211;
  assign dataArray_33_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_14_cachedata_MPORT_en = dataArray_33_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_14_cachedata_MPORT_addr = dataArray_33_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_14_cachedata_MPORT_data = dataArray_33_14[dataArray_33_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_14_MPORT_addr = replace_set;
  assign dataArray_33_14_MPORT_mask = _GEN_8240 & _GEN_7213;
  assign dataArray_33_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_33_15_cachedata_MPORT_en = dataArray_33_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_33_15_cachedata_MPORT_addr = dataArray_33_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_33_15_cachedata_MPORT_data = dataArray_33_15[dataArray_33_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_33_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_33_15_MPORT_addr = replace_set;
  assign dataArray_33_15_MPORT_mask = _GEN_8240 & _GEN_7215;
  assign dataArray_33_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_0_cachedata_MPORT_en = dataArray_34_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_0_cachedata_MPORT_addr = dataArray_34_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_0_cachedata_MPORT_data = dataArray_34_0[dataArray_34_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_0_MPORT_addr = replace_set;
  assign dataArray_34_0_MPORT_mask = _GEN_8272 & _GEN_7185;
  assign dataArray_34_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_1_cachedata_MPORT_en = dataArray_34_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_1_cachedata_MPORT_addr = dataArray_34_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_1_cachedata_MPORT_data = dataArray_34_1[dataArray_34_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_1_MPORT_addr = replace_set;
  assign dataArray_34_1_MPORT_mask = _GEN_8272 & _GEN_7187;
  assign dataArray_34_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_2_cachedata_MPORT_en = dataArray_34_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_2_cachedata_MPORT_addr = dataArray_34_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_2_cachedata_MPORT_data = dataArray_34_2[dataArray_34_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_2_MPORT_addr = replace_set;
  assign dataArray_34_2_MPORT_mask = _GEN_8272 & _GEN_7189;
  assign dataArray_34_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_3_cachedata_MPORT_en = dataArray_34_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_3_cachedata_MPORT_addr = dataArray_34_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_3_cachedata_MPORT_data = dataArray_34_3[dataArray_34_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_3_MPORT_addr = replace_set;
  assign dataArray_34_3_MPORT_mask = _GEN_8272 & _GEN_7191;
  assign dataArray_34_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_4_cachedata_MPORT_en = dataArray_34_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_4_cachedata_MPORT_addr = dataArray_34_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_4_cachedata_MPORT_data = dataArray_34_4[dataArray_34_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_4_MPORT_addr = replace_set;
  assign dataArray_34_4_MPORT_mask = _GEN_8272 & _GEN_7193;
  assign dataArray_34_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_5_cachedata_MPORT_en = dataArray_34_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_5_cachedata_MPORT_addr = dataArray_34_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_5_cachedata_MPORT_data = dataArray_34_5[dataArray_34_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_5_MPORT_addr = replace_set;
  assign dataArray_34_5_MPORT_mask = _GEN_8272 & _GEN_7195;
  assign dataArray_34_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_6_cachedata_MPORT_en = dataArray_34_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_6_cachedata_MPORT_addr = dataArray_34_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_6_cachedata_MPORT_data = dataArray_34_6[dataArray_34_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_6_MPORT_addr = replace_set;
  assign dataArray_34_6_MPORT_mask = _GEN_8272 & _GEN_7197;
  assign dataArray_34_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_7_cachedata_MPORT_en = dataArray_34_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_7_cachedata_MPORT_addr = dataArray_34_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_7_cachedata_MPORT_data = dataArray_34_7[dataArray_34_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_7_MPORT_addr = replace_set;
  assign dataArray_34_7_MPORT_mask = _GEN_8272 & _GEN_7199;
  assign dataArray_34_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_8_cachedata_MPORT_en = dataArray_34_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_8_cachedata_MPORT_addr = dataArray_34_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_8_cachedata_MPORT_data = dataArray_34_8[dataArray_34_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_8_MPORT_addr = replace_set;
  assign dataArray_34_8_MPORT_mask = _GEN_8272 & _GEN_7201;
  assign dataArray_34_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_9_cachedata_MPORT_en = dataArray_34_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_9_cachedata_MPORT_addr = dataArray_34_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_9_cachedata_MPORT_data = dataArray_34_9[dataArray_34_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_9_MPORT_addr = replace_set;
  assign dataArray_34_9_MPORT_mask = _GEN_8272 & _GEN_7203;
  assign dataArray_34_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_10_cachedata_MPORT_en = dataArray_34_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_10_cachedata_MPORT_addr = dataArray_34_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_10_cachedata_MPORT_data = dataArray_34_10[dataArray_34_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_10_MPORT_addr = replace_set;
  assign dataArray_34_10_MPORT_mask = _GEN_8272 & _GEN_7205;
  assign dataArray_34_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_11_cachedata_MPORT_en = dataArray_34_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_11_cachedata_MPORT_addr = dataArray_34_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_11_cachedata_MPORT_data = dataArray_34_11[dataArray_34_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_11_MPORT_addr = replace_set;
  assign dataArray_34_11_MPORT_mask = _GEN_8272 & _GEN_7207;
  assign dataArray_34_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_12_cachedata_MPORT_en = dataArray_34_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_12_cachedata_MPORT_addr = dataArray_34_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_12_cachedata_MPORT_data = dataArray_34_12[dataArray_34_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_12_MPORT_addr = replace_set;
  assign dataArray_34_12_MPORT_mask = _GEN_8272 & _GEN_7209;
  assign dataArray_34_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_13_cachedata_MPORT_en = dataArray_34_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_13_cachedata_MPORT_addr = dataArray_34_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_13_cachedata_MPORT_data = dataArray_34_13[dataArray_34_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_13_MPORT_addr = replace_set;
  assign dataArray_34_13_MPORT_mask = _GEN_8272 & _GEN_7211;
  assign dataArray_34_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_14_cachedata_MPORT_en = dataArray_34_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_14_cachedata_MPORT_addr = dataArray_34_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_14_cachedata_MPORT_data = dataArray_34_14[dataArray_34_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_14_MPORT_addr = replace_set;
  assign dataArray_34_14_MPORT_mask = _GEN_8272 & _GEN_7213;
  assign dataArray_34_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_34_15_cachedata_MPORT_en = dataArray_34_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_34_15_cachedata_MPORT_addr = dataArray_34_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_34_15_cachedata_MPORT_data = dataArray_34_15[dataArray_34_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_34_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_34_15_MPORT_addr = replace_set;
  assign dataArray_34_15_MPORT_mask = _GEN_8272 & _GEN_7215;
  assign dataArray_34_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_0_cachedata_MPORT_en = dataArray_35_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_0_cachedata_MPORT_addr = dataArray_35_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_0_cachedata_MPORT_data = dataArray_35_0[dataArray_35_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_0_MPORT_addr = replace_set;
  assign dataArray_35_0_MPORT_mask = _GEN_8304 & _GEN_7185;
  assign dataArray_35_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_1_cachedata_MPORT_en = dataArray_35_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_1_cachedata_MPORT_addr = dataArray_35_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_1_cachedata_MPORT_data = dataArray_35_1[dataArray_35_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_1_MPORT_addr = replace_set;
  assign dataArray_35_1_MPORT_mask = _GEN_8304 & _GEN_7187;
  assign dataArray_35_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_2_cachedata_MPORT_en = dataArray_35_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_2_cachedata_MPORT_addr = dataArray_35_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_2_cachedata_MPORT_data = dataArray_35_2[dataArray_35_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_2_MPORT_addr = replace_set;
  assign dataArray_35_2_MPORT_mask = _GEN_8304 & _GEN_7189;
  assign dataArray_35_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_3_cachedata_MPORT_en = dataArray_35_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_3_cachedata_MPORT_addr = dataArray_35_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_3_cachedata_MPORT_data = dataArray_35_3[dataArray_35_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_3_MPORT_addr = replace_set;
  assign dataArray_35_3_MPORT_mask = _GEN_8304 & _GEN_7191;
  assign dataArray_35_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_4_cachedata_MPORT_en = dataArray_35_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_4_cachedata_MPORT_addr = dataArray_35_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_4_cachedata_MPORT_data = dataArray_35_4[dataArray_35_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_4_MPORT_addr = replace_set;
  assign dataArray_35_4_MPORT_mask = _GEN_8304 & _GEN_7193;
  assign dataArray_35_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_5_cachedata_MPORT_en = dataArray_35_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_5_cachedata_MPORT_addr = dataArray_35_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_5_cachedata_MPORT_data = dataArray_35_5[dataArray_35_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_5_MPORT_addr = replace_set;
  assign dataArray_35_5_MPORT_mask = _GEN_8304 & _GEN_7195;
  assign dataArray_35_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_6_cachedata_MPORT_en = dataArray_35_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_6_cachedata_MPORT_addr = dataArray_35_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_6_cachedata_MPORT_data = dataArray_35_6[dataArray_35_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_6_MPORT_addr = replace_set;
  assign dataArray_35_6_MPORT_mask = _GEN_8304 & _GEN_7197;
  assign dataArray_35_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_7_cachedata_MPORT_en = dataArray_35_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_7_cachedata_MPORT_addr = dataArray_35_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_7_cachedata_MPORT_data = dataArray_35_7[dataArray_35_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_7_MPORT_addr = replace_set;
  assign dataArray_35_7_MPORT_mask = _GEN_8304 & _GEN_7199;
  assign dataArray_35_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_8_cachedata_MPORT_en = dataArray_35_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_8_cachedata_MPORT_addr = dataArray_35_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_8_cachedata_MPORT_data = dataArray_35_8[dataArray_35_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_8_MPORT_addr = replace_set;
  assign dataArray_35_8_MPORT_mask = _GEN_8304 & _GEN_7201;
  assign dataArray_35_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_9_cachedata_MPORT_en = dataArray_35_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_9_cachedata_MPORT_addr = dataArray_35_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_9_cachedata_MPORT_data = dataArray_35_9[dataArray_35_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_9_MPORT_addr = replace_set;
  assign dataArray_35_9_MPORT_mask = _GEN_8304 & _GEN_7203;
  assign dataArray_35_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_10_cachedata_MPORT_en = dataArray_35_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_10_cachedata_MPORT_addr = dataArray_35_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_10_cachedata_MPORT_data = dataArray_35_10[dataArray_35_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_10_MPORT_addr = replace_set;
  assign dataArray_35_10_MPORT_mask = _GEN_8304 & _GEN_7205;
  assign dataArray_35_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_11_cachedata_MPORT_en = dataArray_35_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_11_cachedata_MPORT_addr = dataArray_35_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_11_cachedata_MPORT_data = dataArray_35_11[dataArray_35_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_11_MPORT_addr = replace_set;
  assign dataArray_35_11_MPORT_mask = _GEN_8304 & _GEN_7207;
  assign dataArray_35_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_12_cachedata_MPORT_en = dataArray_35_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_12_cachedata_MPORT_addr = dataArray_35_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_12_cachedata_MPORT_data = dataArray_35_12[dataArray_35_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_12_MPORT_addr = replace_set;
  assign dataArray_35_12_MPORT_mask = _GEN_8304 & _GEN_7209;
  assign dataArray_35_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_13_cachedata_MPORT_en = dataArray_35_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_13_cachedata_MPORT_addr = dataArray_35_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_13_cachedata_MPORT_data = dataArray_35_13[dataArray_35_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_13_MPORT_addr = replace_set;
  assign dataArray_35_13_MPORT_mask = _GEN_8304 & _GEN_7211;
  assign dataArray_35_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_14_cachedata_MPORT_en = dataArray_35_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_14_cachedata_MPORT_addr = dataArray_35_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_14_cachedata_MPORT_data = dataArray_35_14[dataArray_35_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_14_MPORT_addr = replace_set;
  assign dataArray_35_14_MPORT_mask = _GEN_8304 & _GEN_7213;
  assign dataArray_35_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_35_15_cachedata_MPORT_en = dataArray_35_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_35_15_cachedata_MPORT_addr = dataArray_35_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_35_15_cachedata_MPORT_data = dataArray_35_15[dataArray_35_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_35_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_35_15_MPORT_addr = replace_set;
  assign dataArray_35_15_MPORT_mask = _GEN_8304 & _GEN_7215;
  assign dataArray_35_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_0_cachedata_MPORT_en = dataArray_36_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_0_cachedata_MPORT_addr = dataArray_36_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_0_cachedata_MPORT_data = dataArray_36_0[dataArray_36_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_0_MPORT_addr = replace_set;
  assign dataArray_36_0_MPORT_mask = _GEN_8336 & _GEN_7185;
  assign dataArray_36_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_1_cachedata_MPORT_en = dataArray_36_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_1_cachedata_MPORT_addr = dataArray_36_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_1_cachedata_MPORT_data = dataArray_36_1[dataArray_36_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_1_MPORT_addr = replace_set;
  assign dataArray_36_1_MPORT_mask = _GEN_8336 & _GEN_7187;
  assign dataArray_36_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_2_cachedata_MPORT_en = dataArray_36_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_2_cachedata_MPORT_addr = dataArray_36_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_2_cachedata_MPORT_data = dataArray_36_2[dataArray_36_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_2_MPORT_addr = replace_set;
  assign dataArray_36_2_MPORT_mask = _GEN_8336 & _GEN_7189;
  assign dataArray_36_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_3_cachedata_MPORT_en = dataArray_36_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_3_cachedata_MPORT_addr = dataArray_36_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_3_cachedata_MPORT_data = dataArray_36_3[dataArray_36_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_3_MPORT_addr = replace_set;
  assign dataArray_36_3_MPORT_mask = _GEN_8336 & _GEN_7191;
  assign dataArray_36_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_4_cachedata_MPORT_en = dataArray_36_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_4_cachedata_MPORT_addr = dataArray_36_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_4_cachedata_MPORT_data = dataArray_36_4[dataArray_36_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_4_MPORT_addr = replace_set;
  assign dataArray_36_4_MPORT_mask = _GEN_8336 & _GEN_7193;
  assign dataArray_36_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_5_cachedata_MPORT_en = dataArray_36_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_5_cachedata_MPORT_addr = dataArray_36_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_5_cachedata_MPORT_data = dataArray_36_5[dataArray_36_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_5_MPORT_addr = replace_set;
  assign dataArray_36_5_MPORT_mask = _GEN_8336 & _GEN_7195;
  assign dataArray_36_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_6_cachedata_MPORT_en = dataArray_36_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_6_cachedata_MPORT_addr = dataArray_36_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_6_cachedata_MPORT_data = dataArray_36_6[dataArray_36_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_6_MPORT_addr = replace_set;
  assign dataArray_36_6_MPORT_mask = _GEN_8336 & _GEN_7197;
  assign dataArray_36_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_7_cachedata_MPORT_en = dataArray_36_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_7_cachedata_MPORT_addr = dataArray_36_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_7_cachedata_MPORT_data = dataArray_36_7[dataArray_36_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_7_MPORT_addr = replace_set;
  assign dataArray_36_7_MPORT_mask = _GEN_8336 & _GEN_7199;
  assign dataArray_36_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_8_cachedata_MPORT_en = dataArray_36_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_8_cachedata_MPORT_addr = dataArray_36_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_8_cachedata_MPORT_data = dataArray_36_8[dataArray_36_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_8_MPORT_addr = replace_set;
  assign dataArray_36_8_MPORT_mask = _GEN_8336 & _GEN_7201;
  assign dataArray_36_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_9_cachedata_MPORT_en = dataArray_36_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_9_cachedata_MPORT_addr = dataArray_36_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_9_cachedata_MPORT_data = dataArray_36_9[dataArray_36_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_9_MPORT_addr = replace_set;
  assign dataArray_36_9_MPORT_mask = _GEN_8336 & _GEN_7203;
  assign dataArray_36_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_10_cachedata_MPORT_en = dataArray_36_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_10_cachedata_MPORT_addr = dataArray_36_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_10_cachedata_MPORT_data = dataArray_36_10[dataArray_36_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_10_MPORT_addr = replace_set;
  assign dataArray_36_10_MPORT_mask = _GEN_8336 & _GEN_7205;
  assign dataArray_36_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_11_cachedata_MPORT_en = dataArray_36_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_11_cachedata_MPORT_addr = dataArray_36_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_11_cachedata_MPORT_data = dataArray_36_11[dataArray_36_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_11_MPORT_addr = replace_set;
  assign dataArray_36_11_MPORT_mask = _GEN_8336 & _GEN_7207;
  assign dataArray_36_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_12_cachedata_MPORT_en = dataArray_36_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_12_cachedata_MPORT_addr = dataArray_36_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_12_cachedata_MPORT_data = dataArray_36_12[dataArray_36_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_12_MPORT_addr = replace_set;
  assign dataArray_36_12_MPORT_mask = _GEN_8336 & _GEN_7209;
  assign dataArray_36_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_13_cachedata_MPORT_en = dataArray_36_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_13_cachedata_MPORT_addr = dataArray_36_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_13_cachedata_MPORT_data = dataArray_36_13[dataArray_36_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_13_MPORT_addr = replace_set;
  assign dataArray_36_13_MPORT_mask = _GEN_8336 & _GEN_7211;
  assign dataArray_36_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_14_cachedata_MPORT_en = dataArray_36_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_14_cachedata_MPORT_addr = dataArray_36_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_14_cachedata_MPORT_data = dataArray_36_14[dataArray_36_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_14_MPORT_addr = replace_set;
  assign dataArray_36_14_MPORT_mask = _GEN_8336 & _GEN_7213;
  assign dataArray_36_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_36_15_cachedata_MPORT_en = dataArray_36_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_36_15_cachedata_MPORT_addr = dataArray_36_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_36_15_cachedata_MPORT_data = dataArray_36_15[dataArray_36_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_36_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_36_15_MPORT_addr = replace_set;
  assign dataArray_36_15_MPORT_mask = _GEN_8336 & _GEN_7215;
  assign dataArray_36_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_0_cachedata_MPORT_en = dataArray_37_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_0_cachedata_MPORT_addr = dataArray_37_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_0_cachedata_MPORT_data = dataArray_37_0[dataArray_37_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_0_MPORT_addr = replace_set;
  assign dataArray_37_0_MPORT_mask = _GEN_8368 & _GEN_7185;
  assign dataArray_37_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_1_cachedata_MPORT_en = dataArray_37_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_1_cachedata_MPORT_addr = dataArray_37_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_1_cachedata_MPORT_data = dataArray_37_1[dataArray_37_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_1_MPORT_addr = replace_set;
  assign dataArray_37_1_MPORT_mask = _GEN_8368 & _GEN_7187;
  assign dataArray_37_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_2_cachedata_MPORT_en = dataArray_37_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_2_cachedata_MPORT_addr = dataArray_37_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_2_cachedata_MPORT_data = dataArray_37_2[dataArray_37_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_2_MPORT_addr = replace_set;
  assign dataArray_37_2_MPORT_mask = _GEN_8368 & _GEN_7189;
  assign dataArray_37_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_3_cachedata_MPORT_en = dataArray_37_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_3_cachedata_MPORT_addr = dataArray_37_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_3_cachedata_MPORT_data = dataArray_37_3[dataArray_37_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_3_MPORT_addr = replace_set;
  assign dataArray_37_3_MPORT_mask = _GEN_8368 & _GEN_7191;
  assign dataArray_37_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_4_cachedata_MPORT_en = dataArray_37_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_4_cachedata_MPORT_addr = dataArray_37_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_4_cachedata_MPORT_data = dataArray_37_4[dataArray_37_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_4_MPORT_addr = replace_set;
  assign dataArray_37_4_MPORT_mask = _GEN_8368 & _GEN_7193;
  assign dataArray_37_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_5_cachedata_MPORT_en = dataArray_37_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_5_cachedata_MPORT_addr = dataArray_37_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_5_cachedata_MPORT_data = dataArray_37_5[dataArray_37_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_5_MPORT_addr = replace_set;
  assign dataArray_37_5_MPORT_mask = _GEN_8368 & _GEN_7195;
  assign dataArray_37_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_6_cachedata_MPORT_en = dataArray_37_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_6_cachedata_MPORT_addr = dataArray_37_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_6_cachedata_MPORT_data = dataArray_37_6[dataArray_37_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_6_MPORT_addr = replace_set;
  assign dataArray_37_6_MPORT_mask = _GEN_8368 & _GEN_7197;
  assign dataArray_37_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_7_cachedata_MPORT_en = dataArray_37_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_7_cachedata_MPORT_addr = dataArray_37_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_7_cachedata_MPORT_data = dataArray_37_7[dataArray_37_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_7_MPORT_addr = replace_set;
  assign dataArray_37_7_MPORT_mask = _GEN_8368 & _GEN_7199;
  assign dataArray_37_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_8_cachedata_MPORT_en = dataArray_37_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_8_cachedata_MPORT_addr = dataArray_37_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_8_cachedata_MPORT_data = dataArray_37_8[dataArray_37_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_8_MPORT_addr = replace_set;
  assign dataArray_37_8_MPORT_mask = _GEN_8368 & _GEN_7201;
  assign dataArray_37_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_9_cachedata_MPORT_en = dataArray_37_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_9_cachedata_MPORT_addr = dataArray_37_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_9_cachedata_MPORT_data = dataArray_37_9[dataArray_37_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_9_MPORT_addr = replace_set;
  assign dataArray_37_9_MPORT_mask = _GEN_8368 & _GEN_7203;
  assign dataArray_37_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_10_cachedata_MPORT_en = dataArray_37_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_10_cachedata_MPORT_addr = dataArray_37_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_10_cachedata_MPORT_data = dataArray_37_10[dataArray_37_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_10_MPORT_addr = replace_set;
  assign dataArray_37_10_MPORT_mask = _GEN_8368 & _GEN_7205;
  assign dataArray_37_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_11_cachedata_MPORT_en = dataArray_37_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_11_cachedata_MPORT_addr = dataArray_37_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_11_cachedata_MPORT_data = dataArray_37_11[dataArray_37_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_11_MPORT_addr = replace_set;
  assign dataArray_37_11_MPORT_mask = _GEN_8368 & _GEN_7207;
  assign dataArray_37_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_12_cachedata_MPORT_en = dataArray_37_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_12_cachedata_MPORT_addr = dataArray_37_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_12_cachedata_MPORT_data = dataArray_37_12[dataArray_37_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_12_MPORT_addr = replace_set;
  assign dataArray_37_12_MPORT_mask = _GEN_8368 & _GEN_7209;
  assign dataArray_37_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_13_cachedata_MPORT_en = dataArray_37_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_13_cachedata_MPORT_addr = dataArray_37_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_13_cachedata_MPORT_data = dataArray_37_13[dataArray_37_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_13_MPORT_addr = replace_set;
  assign dataArray_37_13_MPORT_mask = _GEN_8368 & _GEN_7211;
  assign dataArray_37_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_14_cachedata_MPORT_en = dataArray_37_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_14_cachedata_MPORT_addr = dataArray_37_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_14_cachedata_MPORT_data = dataArray_37_14[dataArray_37_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_14_MPORT_addr = replace_set;
  assign dataArray_37_14_MPORT_mask = _GEN_8368 & _GEN_7213;
  assign dataArray_37_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_37_15_cachedata_MPORT_en = dataArray_37_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_37_15_cachedata_MPORT_addr = dataArray_37_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_37_15_cachedata_MPORT_data = dataArray_37_15[dataArray_37_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_37_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_37_15_MPORT_addr = replace_set;
  assign dataArray_37_15_MPORT_mask = _GEN_8368 & _GEN_7215;
  assign dataArray_37_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_0_cachedata_MPORT_en = dataArray_38_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_0_cachedata_MPORT_addr = dataArray_38_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_0_cachedata_MPORT_data = dataArray_38_0[dataArray_38_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_0_MPORT_addr = replace_set;
  assign dataArray_38_0_MPORT_mask = _GEN_8400 & _GEN_7185;
  assign dataArray_38_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_1_cachedata_MPORT_en = dataArray_38_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_1_cachedata_MPORT_addr = dataArray_38_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_1_cachedata_MPORT_data = dataArray_38_1[dataArray_38_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_1_MPORT_addr = replace_set;
  assign dataArray_38_1_MPORT_mask = _GEN_8400 & _GEN_7187;
  assign dataArray_38_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_2_cachedata_MPORT_en = dataArray_38_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_2_cachedata_MPORT_addr = dataArray_38_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_2_cachedata_MPORT_data = dataArray_38_2[dataArray_38_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_2_MPORT_addr = replace_set;
  assign dataArray_38_2_MPORT_mask = _GEN_8400 & _GEN_7189;
  assign dataArray_38_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_3_cachedata_MPORT_en = dataArray_38_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_3_cachedata_MPORT_addr = dataArray_38_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_3_cachedata_MPORT_data = dataArray_38_3[dataArray_38_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_3_MPORT_addr = replace_set;
  assign dataArray_38_3_MPORT_mask = _GEN_8400 & _GEN_7191;
  assign dataArray_38_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_4_cachedata_MPORT_en = dataArray_38_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_4_cachedata_MPORT_addr = dataArray_38_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_4_cachedata_MPORT_data = dataArray_38_4[dataArray_38_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_4_MPORT_addr = replace_set;
  assign dataArray_38_4_MPORT_mask = _GEN_8400 & _GEN_7193;
  assign dataArray_38_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_5_cachedata_MPORT_en = dataArray_38_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_5_cachedata_MPORT_addr = dataArray_38_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_5_cachedata_MPORT_data = dataArray_38_5[dataArray_38_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_5_MPORT_addr = replace_set;
  assign dataArray_38_5_MPORT_mask = _GEN_8400 & _GEN_7195;
  assign dataArray_38_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_6_cachedata_MPORT_en = dataArray_38_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_6_cachedata_MPORT_addr = dataArray_38_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_6_cachedata_MPORT_data = dataArray_38_6[dataArray_38_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_6_MPORT_addr = replace_set;
  assign dataArray_38_6_MPORT_mask = _GEN_8400 & _GEN_7197;
  assign dataArray_38_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_7_cachedata_MPORT_en = dataArray_38_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_7_cachedata_MPORT_addr = dataArray_38_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_7_cachedata_MPORT_data = dataArray_38_7[dataArray_38_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_7_MPORT_addr = replace_set;
  assign dataArray_38_7_MPORT_mask = _GEN_8400 & _GEN_7199;
  assign dataArray_38_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_8_cachedata_MPORT_en = dataArray_38_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_8_cachedata_MPORT_addr = dataArray_38_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_8_cachedata_MPORT_data = dataArray_38_8[dataArray_38_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_8_MPORT_addr = replace_set;
  assign dataArray_38_8_MPORT_mask = _GEN_8400 & _GEN_7201;
  assign dataArray_38_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_9_cachedata_MPORT_en = dataArray_38_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_9_cachedata_MPORT_addr = dataArray_38_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_9_cachedata_MPORT_data = dataArray_38_9[dataArray_38_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_9_MPORT_addr = replace_set;
  assign dataArray_38_9_MPORT_mask = _GEN_8400 & _GEN_7203;
  assign dataArray_38_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_10_cachedata_MPORT_en = dataArray_38_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_10_cachedata_MPORT_addr = dataArray_38_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_10_cachedata_MPORT_data = dataArray_38_10[dataArray_38_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_10_MPORT_addr = replace_set;
  assign dataArray_38_10_MPORT_mask = _GEN_8400 & _GEN_7205;
  assign dataArray_38_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_11_cachedata_MPORT_en = dataArray_38_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_11_cachedata_MPORT_addr = dataArray_38_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_11_cachedata_MPORT_data = dataArray_38_11[dataArray_38_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_11_MPORT_addr = replace_set;
  assign dataArray_38_11_MPORT_mask = _GEN_8400 & _GEN_7207;
  assign dataArray_38_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_12_cachedata_MPORT_en = dataArray_38_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_12_cachedata_MPORT_addr = dataArray_38_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_12_cachedata_MPORT_data = dataArray_38_12[dataArray_38_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_12_MPORT_addr = replace_set;
  assign dataArray_38_12_MPORT_mask = _GEN_8400 & _GEN_7209;
  assign dataArray_38_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_13_cachedata_MPORT_en = dataArray_38_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_13_cachedata_MPORT_addr = dataArray_38_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_13_cachedata_MPORT_data = dataArray_38_13[dataArray_38_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_13_MPORT_addr = replace_set;
  assign dataArray_38_13_MPORT_mask = _GEN_8400 & _GEN_7211;
  assign dataArray_38_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_14_cachedata_MPORT_en = dataArray_38_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_14_cachedata_MPORT_addr = dataArray_38_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_14_cachedata_MPORT_data = dataArray_38_14[dataArray_38_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_14_MPORT_addr = replace_set;
  assign dataArray_38_14_MPORT_mask = _GEN_8400 & _GEN_7213;
  assign dataArray_38_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_38_15_cachedata_MPORT_en = dataArray_38_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_38_15_cachedata_MPORT_addr = dataArray_38_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_38_15_cachedata_MPORT_data = dataArray_38_15[dataArray_38_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_38_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_38_15_MPORT_addr = replace_set;
  assign dataArray_38_15_MPORT_mask = _GEN_8400 & _GEN_7215;
  assign dataArray_38_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_0_cachedata_MPORT_en = dataArray_39_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_0_cachedata_MPORT_addr = dataArray_39_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_0_cachedata_MPORT_data = dataArray_39_0[dataArray_39_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_0_MPORT_addr = replace_set;
  assign dataArray_39_0_MPORT_mask = _GEN_8432 & _GEN_7185;
  assign dataArray_39_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_1_cachedata_MPORT_en = dataArray_39_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_1_cachedata_MPORT_addr = dataArray_39_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_1_cachedata_MPORT_data = dataArray_39_1[dataArray_39_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_1_MPORT_addr = replace_set;
  assign dataArray_39_1_MPORT_mask = _GEN_8432 & _GEN_7187;
  assign dataArray_39_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_2_cachedata_MPORT_en = dataArray_39_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_2_cachedata_MPORT_addr = dataArray_39_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_2_cachedata_MPORT_data = dataArray_39_2[dataArray_39_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_2_MPORT_addr = replace_set;
  assign dataArray_39_2_MPORT_mask = _GEN_8432 & _GEN_7189;
  assign dataArray_39_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_3_cachedata_MPORT_en = dataArray_39_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_3_cachedata_MPORT_addr = dataArray_39_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_3_cachedata_MPORT_data = dataArray_39_3[dataArray_39_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_3_MPORT_addr = replace_set;
  assign dataArray_39_3_MPORT_mask = _GEN_8432 & _GEN_7191;
  assign dataArray_39_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_4_cachedata_MPORT_en = dataArray_39_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_4_cachedata_MPORT_addr = dataArray_39_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_4_cachedata_MPORT_data = dataArray_39_4[dataArray_39_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_4_MPORT_addr = replace_set;
  assign dataArray_39_4_MPORT_mask = _GEN_8432 & _GEN_7193;
  assign dataArray_39_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_5_cachedata_MPORT_en = dataArray_39_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_5_cachedata_MPORT_addr = dataArray_39_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_5_cachedata_MPORT_data = dataArray_39_5[dataArray_39_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_5_MPORT_addr = replace_set;
  assign dataArray_39_5_MPORT_mask = _GEN_8432 & _GEN_7195;
  assign dataArray_39_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_6_cachedata_MPORT_en = dataArray_39_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_6_cachedata_MPORT_addr = dataArray_39_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_6_cachedata_MPORT_data = dataArray_39_6[dataArray_39_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_6_MPORT_addr = replace_set;
  assign dataArray_39_6_MPORT_mask = _GEN_8432 & _GEN_7197;
  assign dataArray_39_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_7_cachedata_MPORT_en = dataArray_39_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_7_cachedata_MPORT_addr = dataArray_39_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_7_cachedata_MPORT_data = dataArray_39_7[dataArray_39_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_7_MPORT_addr = replace_set;
  assign dataArray_39_7_MPORT_mask = _GEN_8432 & _GEN_7199;
  assign dataArray_39_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_8_cachedata_MPORT_en = dataArray_39_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_8_cachedata_MPORT_addr = dataArray_39_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_8_cachedata_MPORT_data = dataArray_39_8[dataArray_39_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_8_MPORT_addr = replace_set;
  assign dataArray_39_8_MPORT_mask = _GEN_8432 & _GEN_7201;
  assign dataArray_39_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_9_cachedata_MPORT_en = dataArray_39_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_9_cachedata_MPORT_addr = dataArray_39_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_9_cachedata_MPORT_data = dataArray_39_9[dataArray_39_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_9_MPORT_addr = replace_set;
  assign dataArray_39_9_MPORT_mask = _GEN_8432 & _GEN_7203;
  assign dataArray_39_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_10_cachedata_MPORT_en = dataArray_39_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_10_cachedata_MPORT_addr = dataArray_39_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_10_cachedata_MPORT_data = dataArray_39_10[dataArray_39_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_10_MPORT_addr = replace_set;
  assign dataArray_39_10_MPORT_mask = _GEN_8432 & _GEN_7205;
  assign dataArray_39_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_11_cachedata_MPORT_en = dataArray_39_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_11_cachedata_MPORT_addr = dataArray_39_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_11_cachedata_MPORT_data = dataArray_39_11[dataArray_39_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_11_MPORT_addr = replace_set;
  assign dataArray_39_11_MPORT_mask = _GEN_8432 & _GEN_7207;
  assign dataArray_39_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_12_cachedata_MPORT_en = dataArray_39_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_12_cachedata_MPORT_addr = dataArray_39_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_12_cachedata_MPORT_data = dataArray_39_12[dataArray_39_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_12_MPORT_addr = replace_set;
  assign dataArray_39_12_MPORT_mask = _GEN_8432 & _GEN_7209;
  assign dataArray_39_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_13_cachedata_MPORT_en = dataArray_39_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_13_cachedata_MPORT_addr = dataArray_39_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_13_cachedata_MPORT_data = dataArray_39_13[dataArray_39_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_13_MPORT_addr = replace_set;
  assign dataArray_39_13_MPORT_mask = _GEN_8432 & _GEN_7211;
  assign dataArray_39_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_14_cachedata_MPORT_en = dataArray_39_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_14_cachedata_MPORT_addr = dataArray_39_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_14_cachedata_MPORT_data = dataArray_39_14[dataArray_39_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_14_MPORT_addr = replace_set;
  assign dataArray_39_14_MPORT_mask = _GEN_8432 & _GEN_7213;
  assign dataArray_39_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_39_15_cachedata_MPORT_en = dataArray_39_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_39_15_cachedata_MPORT_addr = dataArray_39_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_39_15_cachedata_MPORT_data = dataArray_39_15[dataArray_39_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_39_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_39_15_MPORT_addr = replace_set;
  assign dataArray_39_15_MPORT_mask = _GEN_8432 & _GEN_7215;
  assign dataArray_39_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_0_cachedata_MPORT_en = dataArray_40_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_0_cachedata_MPORT_addr = dataArray_40_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_0_cachedata_MPORT_data = dataArray_40_0[dataArray_40_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_0_MPORT_addr = replace_set;
  assign dataArray_40_0_MPORT_mask = _GEN_8464 & _GEN_7185;
  assign dataArray_40_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_1_cachedata_MPORT_en = dataArray_40_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_1_cachedata_MPORT_addr = dataArray_40_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_1_cachedata_MPORT_data = dataArray_40_1[dataArray_40_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_1_MPORT_addr = replace_set;
  assign dataArray_40_1_MPORT_mask = _GEN_8464 & _GEN_7187;
  assign dataArray_40_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_2_cachedata_MPORT_en = dataArray_40_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_2_cachedata_MPORT_addr = dataArray_40_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_2_cachedata_MPORT_data = dataArray_40_2[dataArray_40_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_2_MPORT_addr = replace_set;
  assign dataArray_40_2_MPORT_mask = _GEN_8464 & _GEN_7189;
  assign dataArray_40_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_3_cachedata_MPORT_en = dataArray_40_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_3_cachedata_MPORT_addr = dataArray_40_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_3_cachedata_MPORT_data = dataArray_40_3[dataArray_40_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_3_MPORT_addr = replace_set;
  assign dataArray_40_3_MPORT_mask = _GEN_8464 & _GEN_7191;
  assign dataArray_40_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_4_cachedata_MPORT_en = dataArray_40_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_4_cachedata_MPORT_addr = dataArray_40_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_4_cachedata_MPORT_data = dataArray_40_4[dataArray_40_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_4_MPORT_addr = replace_set;
  assign dataArray_40_4_MPORT_mask = _GEN_8464 & _GEN_7193;
  assign dataArray_40_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_5_cachedata_MPORT_en = dataArray_40_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_5_cachedata_MPORT_addr = dataArray_40_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_5_cachedata_MPORT_data = dataArray_40_5[dataArray_40_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_5_MPORT_addr = replace_set;
  assign dataArray_40_5_MPORT_mask = _GEN_8464 & _GEN_7195;
  assign dataArray_40_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_6_cachedata_MPORT_en = dataArray_40_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_6_cachedata_MPORT_addr = dataArray_40_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_6_cachedata_MPORT_data = dataArray_40_6[dataArray_40_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_6_MPORT_addr = replace_set;
  assign dataArray_40_6_MPORT_mask = _GEN_8464 & _GEN_7197;
  assign dataArray_40_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_7_cachedata_MPORT_en = dataArray_40_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_7_cachedata_MPORT_addr = dataArray_40_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_7_cachedata_MPORT_data = dataArray_40_7[dataArray_40_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_7_MPORT_addr = replace_set;
  assign dataArray_40_7_MPORT_mask = _GEN_8464 & _GEN_7199;
  assign dataArray_40_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_8_cachedata_MPORT_en = dataArray_40_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_8_cachedata_MPORT_addr = dataArray_40_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_8_cachedata_MPORT_data = dataArray_40_8[dataArray_40_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_8_MPORT_addr = replace_set;
  assign dataArray_40_8_MPORT_mask = _GEN_8464 & _GEN_7201;
  assign dataArray_40_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_9_cachedata_MPORT_en = dataArray_40_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_9_cachedata_MPORT_addr = dataArray_40_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_9_cachedata_MPORT_data = dataArray_40_9[dataArray_40_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_9_MPORT_addr = replace_set;
  assign dataArray_40_9_MPORT_mask = _GEN_8464 & _GEN_7203;
  assign dataArray_40_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_10_cachedata_MPORT_en = dataArray_40_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_10_cachedata_MPORT_addr = dataArray_40_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_10_cachedata_MPORT_data = dataArray_40_10[dataArray_40_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_10_MPORT_addr = replace_set;
  assign dataArray_40_10_MPORT_mask = _GEN_8464 & _GEN_7205;
  assign dataArray_40_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_11_cachedata_MPORT_en = dataArray_40_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_11_cachedata_MPORT_addr = dataArray_40_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_11_cachedata_MPORT_data = dataArray_40_11[dataArray_40_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_11_MPORT_addr = replace_set;
  assign dataArray_40_11_MPORT_mask = _GEN_8464 & _GEN_7207;
  assign dataArray_40_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_12_cachedata_MPORT_en = dataArray_40_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_12_cachedata_MPORT_addr = dataArray_40_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_12_cachedata_MPORT_data = dataArray_40_12[dataArray_40_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_12_MPORT_addr = replace_set;
  assign dataArray_40_12_MPORT_mask = _GEN_8464 & _GEN_7209;
  assign dataArray_40_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_13_cachedata_MPORT_en = dataArray_40_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_13_cachedata_MPORT_addr = dataArray_40_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_13_cachedata_MPORT_data = dataArray_40_13[dataArray_40_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_13_MPORT_addr = replace_set;
  assign dataArray_40_13_MPORT_mask = _GEN_8464 & _GEN_7211;
  assign dataArray_40_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_14_cachedata_MPORT_en = dataArray_40_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_14_cachedata_MPORT_addr = dataArray_40_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_14_cachedata_MPORT_data = dataArray_40_14[dataArray_40_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_14_MPORT_addr = replace_set;
  assign dataArray_40_14_MPORT_mask = _GEN_8464 & _GEN_7213;
  assign dataArray_40_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_40_15_cachedata_MPORT_en = dataArray_40_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_40_15_cachedata_MPORT_addr = dataArray_40_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_40_15_cachedata_MPORT_data = dataArray_40_15[dataArray_40_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_40_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_40_15_MPORT_addr = replace_set;
  assign dataArray_40_15_MPORT_mask = _GEN_8464 & _GEN_7215;
  assign dataArray_40_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_0_cachedata_MPORT_en = dataArray_41_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_0_cachedata_MPORT_addr = dataArray_41_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_0_cachedata_MPORT_data = dataArray_41_0[dataArray_41_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_0_MPORT_addr = replace_set;
  assign dataArray_41_0_MPORT_mask = _GEN_8496 & _GEN_7185;
  assign dataArray_41_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_1_cachedata_MPORT_en = dataArray_41_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_1_cachedata_MPORT_addr = dataArray_41_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_1_cachedata_MPORT_data = dataArray_41_1[dataArray_41_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_1_MPORT_addr = replace_set;
  assign dataArray_41_1_MPORT_mask = _GEN_8496 & _GEN_7187;
  assign dataArray_41_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_2_cachedata_MPORT_en = dataArray_41_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_2_cachedata_MPORT_addr = dataArray_41_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_2_cachedata_MPORT_data = dataArray_41_2[dataArray_41_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_2_MPORT_addr = replace_set;
  assign dataArray_41_2_MPORT_mask = _GEN_8496 & _GEN_7189;
  assign dataArray_41_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_3_cachedata_MPORT_en = dataArray_41_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_3_cachedata_MPORT_addr = dataArray_41_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_3_cachedata_MPORT_data = dataArray_41_3[dataArray_41_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_3_MPORT_addr = replace_set;
  assign dataArray_41_3_MPORT_mask = _GEN_8496 & _GEN_7191;
  assign dataArray_41_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_4_cachedata_MPORT_en = dataArray_41_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_4_cachedata_MPORT_addr = dataArray_41_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_4_cachedata_MPORT_data = dataArray_41_4[dataArray_41_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_4_MPORT_addr = replace_set;
  assign dataArray_41_4_MPORT_mask = _GEN_8496 & _GEN_7193;
  assign dataArray_41_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_5_cachedata_MPORT_en = dataArray_41_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_5_cachedata_MPORT_addr = dataArray_41_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_5_cachedata_MPORT_data = dataArray_41_5[dataArray_41_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_5_MPORT_addr = replace_set;
  assign dataArray_41_5_MPORT_mask = _GEN_8496 & _GEN_7195;
  assign dataArray_41_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_6_cachedata_MPORT_en = dataArray_41_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_6_cachedata_MPORT_addr = dataArray_41_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_6_cachedata_MPORT_data = dataArray_41_6[dataArray_41_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_6_MPORT_addr = replace_set;
  assign dataArray_41_6_MPORT_mask = _GEN_8496 & _GEN_7197;
  assign dataArray_41_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_7_cachedata_MPORT_en = dataArray_41_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_7_cachedata_MPORT_addr = dataArray_41_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_7_cachedata_MPORT_data = dataArray_41_7[dataArray_41_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_7_MPORT_addr = replace_set;
  assign dataArray_41_7_MPORT_mask = _GEN_8496 & _GEN_7199;
  assign dataArray_41_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_8_cachedata_MPORT_en = dataArray_41_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_8_cachedata_MPORT_addr = dataArray_41_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_8_cachedata_MPORT_data = dataArray_41_8[dataArray_41_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_8_MPORT_addr = replace_set;
  assign dataArray_41_8_MPORT_mask = _GEN_8496 & _GEN_7201;
  assign dataArray_41_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_9_cachedata_MPORT_en = dataArray_41_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_9_cachedata_MPORT_addr = dataArray_41_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_9_cachedata_MPORT_data = dataArray_41_9[dataArray_41_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_9_MPORT_addr = replace_set;
  assign dataArray_41_9_MPORT_mask = _GEN_8496 & _GEN_7203;
  assign dataArray_41_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_10_cachedata_MPORT_en = dataArray_41_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_10_cachedata_MPORT_addr = dataArray_41_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_10_cachedata_MPORT_data = dataArray_41_10[dataArray_41_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_10_MPORT_addr = replace_set;
  assign dataArray_41_10_MPORT_mask = _GEN_8496 & _GEN_7205;
  assign dataArray_41_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_11_cachedata_MPORT_en = dataArray_41_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_11_cachedata_MPORT_addr = dataArray_41_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_11_cachedata_MPORT_data = dataArray_41_11[dataArray_41_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_11_MPORT_addr = replace_set;
  assign dataArray_41_11_MPORT_mask = _GEN_8496 & _GEN_7207;
  assign dataArray_41_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_12_cachedata_MPORT_en = dataArray_41_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_12_cachedata_MPORT_addr = dataArray_41_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_12_cachedata_MPORT_data = dataArray_41_12[dataArray_41_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_12_MPORT_addr = replace_set;
  assign dataArray_41_12_MPORT_mask = _GEN_8496 & _GEN_7209;
  assign dataArray_41_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_13_cachedata_MPORT_en = dataArray_41_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_13_cachedata_MPORT_addr = dataArray_41_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_13_cachedata_MPORT_data = dataArray_41_13[dataArray_41_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_13_MPORT_addr = replace_set;
  assign dataArray_41_13_MPORT_mask = _GEN_8496 & _GEN_7211;
  assign dataArray_41_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_14_cachedata_MPORT_en = dataArray_41_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_14_cachedata_MPORT_addr = dataArray_41_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_14_cachedata_MPORT_data = dataArray_41_14[dataArray_41_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_14_MPORT_addr = replace_set;
  assign dataArray_41_14_MPORT_mask = _GEN_8496 & _GEN_7213;
  assign dataArray_41_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_41_15_cachedata_MPORT_en = dataArray_41_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_41_15_cachedata_MPORT_addr = dataArray_41_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_41_15_cachedata_MPORT_data = dataArray_41_15[dataArray_41_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_41_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_41_15_MPORT_addr = replace_set;
  assign dataArray_41_15_MPORT_mask = _GEN_8496 & _GEN_7215;
  assign dataArray_41_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_0_cachedata_MPORT_en = dataArray_42_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_0_cachedata_MPORT_addr = dataArray_42_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_0_cachedata_MPORT_data = dataArray_42_0[dataArray_42_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_0_MPORT_addr = replace_set;
  assign dataArray_42_0_MPORT_mask = _GEN_8528 & _GEN_7185;
  assign dataArray_42_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_1_cachedata_MPORT_en = dataArray_42_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_1_cachedata_MPORT_addr = dataArray_42_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_1_cachedata_MPORT_data = dataArray_42_1[dataArray_42_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_1_MPORT_addr = replace_set;
  assign dataArray_42_1_MPORT_mask = _GEN_8528 & _GEN_7187;
  assign dataArray_42_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_2_cachedata_MPORT_en = dataArray_42_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_2_cachedata_MPORT_addr = dataArray_42_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_2_cachedata_MPORT_data = dataArray_42_2[dataArray_42_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_2_MPORT_addr = replace_set;
  assign dataArray_42_2_MPORT_mask = _GEN_8528 & _GEN_7189;
  assign dataArray_42_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_3_cachedata_MPORT_en = dataArray_42_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_3_cachedata_MPORT_addr = dataArray_42_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_3_cachedata_MPORT_data = dataArray_42_3[dataArray_42_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_3_MPORT_addr = replace_set;
  assign dataArray_42_3_MPORT_mask = _GEN_8528 & _GEN_7191;
  assign dataArray_42_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_4_cachedata_MPORT_en = dataArray_42_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_4_cachedata_MPORT_addr = dataArray_42_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_4_cachedata_MPORT_data = dataArray_42_4[dataArray_42_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_4_MPORT_addr = replace_set;
  assign dataArray_42_4_MPORT_mask = _GEN_8528 & _GEN_7193;
  assign dataArray_42_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_5_cachedata_MPORT_en = dataArray_42_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_5_cachedata_MPORT_addr = dataArray_42_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_5_cachedata_MPORT_data = dataArray_42_5[dataArray_42_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_5_MPORT_addr = replace_set;
  assign dataArray_42_5_MPORT_mask = _GEN_8528 & _GEN_7195;
  assign dataArray_42_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_6_cachedata_MPORT_en = dataArray_42_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_6_cachedata_MPORT_addr = dataArray_42_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_6_cachedata_MPORT_data = dataArray_42_6[dataArray_42_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_6_MPORT_addr = replace_set;
  assign dataArray_42_6_MPORT_mask = _GEN_8528 & _GEN_7197;
  assign dataArray_42_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_7_cachedata_MPORT_en = dataArray_42_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_7_cachedata_MPORT_addr = dataArray_42_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_7_cachedata_MPORT_data = dataArray_42_7[dataArray_42_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_7_MPORT_addr = replace_set;
  assign dataArray_42_7_MPORT_mask = _GEN_8528 & _GEN_7199;
  assign dataArray_42_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_8_cachedata_MPORT_en = dataArray_42_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_8_cachedata_MPORT_addr = dataArray_42_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_8_cachedata_MPORT_data = dataArray_42_8[dataArray_42_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_8_MPORT_addr = replace_set;
  assign dataArray_42_8_MPORT_mask = _GEN_8528 & _GEN_7201;
  assign dataArray_42_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_9_cachedata_MPORT_en = dataArray_42_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_9_cachedata_MPORT_addr = dataArray_42_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_9_cachedata_MPORT_data = dataArray_42_9[dataArray_42_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_9_MPORT_addr = replace_set;
  assign dataArray_42_9_MPORT_mask = _GEN_8528 & _GEN_7203;
  assign dataArray_42_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_10_cachedata_MPORT_en = dataArray_42_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_10_cachedata_MPORT_addr = dataArray_42_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_10_cachedata_MPORT_data = dataArray_42_10[dataArray_42_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_10_MPORT_addr = replace_set;
  assign dataArray_42_10_MPORT_mask = _GEN_8528 & _GEN_7205;
  assign dataArray_42_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_11_cachedata_MPORT_en = dataArray_42_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_11_cachedata_MPORT_addr = dataArray_42_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_11_cachedata_MPORT_data = dataArray_42_11[dataArray_42_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_11_MPORT_addr = replace_set;
  assign dataArray_42_11_MPORT_mask = _GEN_8528 & _GEN_7207;
  assign dataArray_42_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_12_cachedata_MPORT_en = dataArray_42_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_12_cachedata_MPORT_addr = dataArray_42_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_12_cachedata_MPORT_data = dataArray_42_12[dataArray_42_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_12_MPORT_addr = replace_set;
  assign dataArray_42_12_MPORT_mask = _GEN_8528 & _GEN_7209;
  assign dataArray_42_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_13_cachedata_MPORT_en = dataArray_42_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_13_cachedata_MPORT_addr = dataArray_42_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_13_cachedata_MPORT_data = dataArray_42_13[dataArray_42_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_13_MPORT_addr = replace_set;
  assign dataArray_42_13_MPORT_mask = _GEN_8528 & _GEN_7211;
  assign dataArray_42_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_14_cachedata_MPORT_en = dataArray_42_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_14_cachedata_MPORT_addr = dataArray_42_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_14_cachedata_MPORT_data = dataArray_42_14[dataArray_42_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_14_MPORT_addr = replace_set;
  assign dataArray_42_14_MPORT_mask = _GEN_8528 & _GEN_7213;
  assign dataArray_42_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_42_15_cachedata_MPORT_en = dataArray_42_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_42_15_cachedata_MPORT_addr = dataArray_42_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_42_15_cachedata_MPORT_data = dataArray_42_15[dataArray_42_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_42_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_42_15_MPORT_addr = replace_set;
  assign dataArray_42_15_MPORT_mask = _GEN_8528 & _GEN_7215;
  assign dataArray_42_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_0_cachedata_MPORT_en = dataArray_43_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_0_cachedata_MPORT_addr = dataArray_43_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_0_cachedata_MPORT_data = dataArray_43_0[dataArray_43_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_0_MPORT_addr = replace_set;
  assign dataArray_43_0_MPORT_mask = _GEN_8560 & _GEN_7185;
  assign dataArray_43_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_1_cachedata_MPORT_en = dataArray_43_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_1_cachedata_MPORT_addr = dataArray_43_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_1_cachedata_MPORT_data = dataArray_43_1[dataArray_43_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_1_MPORT_addr = replace_set;
  assign dataArray_43_1_MPORT_mask = _GEN_8560 & _GEN_7187;
  assign dataArray_43_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_2_cachedata_MPORT_en = dataArray_43_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_2_cachedata_MPORT_addr = dataArray_43_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_2_cachedata_MPORT_data = dataArray_43_2[dataArray_43_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_2_MPORT_addr = replace_set;
  assign dataArray_43_2_MPORT_mask = _GEN_8560 & _GEN_7189;
  assign dataArray_43_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_3_cachedata_MPORT_en = dataArray_43_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_3_cachedata_MPORT_addr = dataArray_43_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_3_cachedata_MPORT_data = dataArray_43_3[dataArray_43_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_3_MPORT_addr = replace_set;
  assign dataArray_43_3_MPORT_mask = _GEN_8560 & _GEN_7191;
  assign dataArray_43_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_4_cachedata_MPORT_en = dataArray_43_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_4_cachedata_MPORT_addr = dataArray_43_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_4_cachedata_MPORT_data = dataArray_43_4[dataArray_43_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_4_MPORT_addr = replace_set;
  assign dataArray_43_4_MPORT_mask = _GEN_8560 & _GEN_7193;
  assign dataArray_43_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_5_cachedata_MPORT_en = dataArray_43_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_5_cachedata_MPORT_addr = dataArray_43_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_5_cachedata_MPORT_data = dataArray_43_5[dataArray_43_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_5_MPORT_addr = replace_set;
  assign dataArray_43_5_MPORT_mask = _GEN_8560 & _GEN_7195;
  assign dataArray_43_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_6_cachedata_MPORT_en = dataArray_43_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_6_cachedata_MPORT_addr = dataArray_43_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_6_cachedata_MPORT_data = dataArray_43_6[dataArray_43_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_6_MPORT_addr = replace_set;
  assign dataArray_43_6_MPORT_mask = _GEN_8560 & _GEN_7197;
  assign dataArray_43_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_7_cachedata_MPORT_en = dataArray_43_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_7_cachedata_MPORT_addr = dataArray_43_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_7_cachedata_MPORT_data = dataArray_43_7[dataArray_43_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_7_MPORT_addr = replace_set;
  assign dataArray_43_7_MPORT_mask = _GEN_8560 & _GEN_7199;
  assign dataArray_43_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_8_cachedata_MPORT_en = dataArray_43_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_8_cachedata_MPORT_addr = dataArray_43_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_8_cachedata_MPORT_data = dataArray_43_8[dataArray_43_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_8_MPORT_addr = replace_set;
  assign dataArray_43_8_MPORT_mask = _GEN_8560 & _GEN_7201;
  assign dataArray_43_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_9_cachedata_MPORT_en = dataArray_43_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_9_cachedata_MPORT_addr = dataArray_43_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_9_cachedata_MPORT_data = dataArray_43_9[dataArray_43_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_9_MPORT_addr = replace_set;
  assign dataArray_43_9_MPORT_mask = _GEN_8560 & _GEN_7203;
  assign dataArray_43_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_10_cachedata_MPORT_en = dataArray_43_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_10_cachedata_MPORT_addr = dataArray_43_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_10_cachedata_MPORT_data = dataArray_43_10[dataArray_43_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_10_MPORT_addr = replace_set;
  assign dataArray_43_10_MPORT_mask = _GEN_8560 & _GEN_7205;
  assign dataArray_43_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_11_cachedata_MPORT_en = dataArray_43_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_11_cachedata_MPORT_addr = dataArray_43_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_11_cachedata_MPORT_data = dataArray_43_11[dataArray_43_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_11_MPORT_addr = replace_set;
  assign dataArray_43_11_MPORT_mask = _GEN_8560 & _GEN_7207;
  assign dataArray_43_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_12_cachedata_MPORT_en = dataArray_43_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_12_cachedata_MPORT_addr = dataArray_43_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_12_cachedata_MPORT_data = dataArray_43_12[dataArray_43_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_12_MPORT_addr = replace_set;
  assign dataArray_43_12_MPORT_mask = _GEN_8560 & _GEN_7209;
  assign dataArray_43_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_13_cachedata_MPORT_en = dataArray_43_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_13_cachedata_MPORT_addr = dataArray_43_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_13_cachedata_MPORT_data = dataArray_43_13[dataArray_43_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_13_MPORT_addr = replace_set;
  assign dataArray_43_13_MPORT_mask = _GEN_8560 & _GEN_7211;
  assign dataArray_43_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_14_cachedata_MPORT_en = dataArray_43_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_14_cachedata_MPORT_addr = dataArray_43_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_14_cachedata_MPORT_data = dataArray_43_14[dataArray_43_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_14_MPORT_addr = replace_set;
  assign dataArray_43_14_MPORT_mask = _GEN_8560 & _GEN_7213;
  assign dataArray_43_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_43_15_cachedata_MPORT_en = dataArray_43_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_43_15_cachedata_MPORT_addr = dataArray_43_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_43_15_cachedata_MPORT_data = dataArray_43_15[dataArray_43_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_43_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_43_15_MPORT_addr = replace_set;
  assign dataArray_43_15_MPORT_mask = _GEN_8560 & _GEN_7215;
  assign dataArray_43_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_0_cachedata_MPORT_en = dataArray_44_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_0_cachedata_MPORT_addr = dataArray_44_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_0_cachedata_MPORT_data = dataArray_44_0[dataArray_44_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_0_MPORT_addr = replace_set;
  assign dataArray_44_0_MPORT_mask = _GEN_8592 & _GEN_7185;
  assign dataArray_44_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_1_cachedata_MPORT_en = dataArray_44_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_1_cachedata_MPORT_addr = dataArray_44_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_1_cachedata_MPORT_data = dataArray_44_1[dataArray_44_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_1_MPORT_addr = replace_set;
  assign dataArray_44_1_MPORT_mask = _GEN_8592 & _GEN_7187;
  assign dataArray_44_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_2_cachedata_MPORT_en = dataArray_44_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_2_cachedata_MPORT_addr = dataArray_44_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_2_cachedata_MPORT_data = dataArray_44_2[dataArray_44_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_2_MPORT_addr = replace_set;
  assign dataArray_44_2_MPORT_mask = _GEN_8592 & _GEN_7189;
  assign dataArray_44_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_3_cachedata_MPORT_en = dataArray_44_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_3_cachedata_MPORT_addr = dataArray_44_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_3_cachedata_MPORT_data = dataArray_44_3[dataArray_44_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_3_MPORT_addr = replace_set;
  assign dataArray_44_3_MPORT_mask = _GEN_8592 & _GEN_7191;
  assign dataArray_44_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_4_cachedata_MPORT_en = dataArray_44_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_4_cachedata_MPORT_addr = dataArray_44_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_4_cachedata_MPORT_data = dataArray_44_4[dataArray_44_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_4_MPORT_addr = replace_set;
  assign dataArray_44_4_MPORT_mask = _GEN_8592 & _GEN_7193;
  assign dataArray_44_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_5_cachedata_MPORT_en = dataArray_44_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_5_cachedata_MPORT_addr = dataArray_44_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_5_cachedata_MPORT_data = dataArray_44_5[dataArray_44_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_5_MPORT_addr = replace_set;
  assign dataArray_44_5_MPORT_mask = _GEN_8592 & _GEN_7195;
  assign dataArray_44_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_6_cachedata_MPORT_en = dataArray_44_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_6_cachedata_MPORT_addr = dataArray_44_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_6_cachedata_MPORT_data = dataArray_44_6[dataArray_44_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_6_MPORT_addr = replace_set;
  assign dataArray_44_6_MPORT_mask = _GEN_8592 & _GEN_7197;
  assign dataArray_44_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_7_cachedata_MPORT_en = dataArray_44_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_7_cachedata_MPORT_addr = dataArray_44_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_7_cachedata_MPORT_data = dataArray_44_7[dataArray_44_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_7_MPORT_addr = replace_set;
  assign dataArray_44_7_MPORT_mask = _GEN_8592 & _GEN_7199;
  assign dataArray_44_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_8_cachedata_MPORT_en = dataArray_44_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_8_cachedata_MPORT_addr = dataArray_44_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_8_cachedata_MPORT_data = dataArray_44_8[dataArray_44_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_8_MPORT_addr = replace_set;
  assign dataArray_44_8_MPORT_mask = _GEN_8592 & _GEN_7201;
  assign dataArray_44_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_9_cachedata_MPORT_en = dataArray_44_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_9_cachedata_MPORT_addr = dataArray_44_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_9_cachedata_MPORT_data = dataArray_44_9[dataArray_44_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_9_MPORT_addr = replace_set;
  assign dataArray_44_9_MPORT_mask = _GEN_8592 & _GEN_7203;
  assign dataArray_44_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_10_cachedata_MPORT_en = dataArray_44_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_10_cachedata_MPORT_addr = dataArray_44_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_10_cachedata_MPORT_data = dataArray_44_10[dataArray_44_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_10_MPORT_addr = replace_set;
  assign dataArray_44_10_MPORT_mask = _GEN_8592 & _GEN_7205;
  assign dataArray_44_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_11_cachedata_MPORT_en = dataArray_44_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_11_cachedata_MPORT_addr = dataArray_44_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_11_cachedata_MPORT_data = dataArray_44_11[dataArray_44_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_11_MPORT_addr = replace_set;
  assign dataArray_44_11_MPORT_mask = _GEN_8592 & _GEN_7207;
  assign dataArray_44_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_12_cachedata_MPORT_en = dataArray_44_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_12_cachedata_MPORT_addr = dataArray_44_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_12_cachedata_MPORT_data = dataArray_44_12[dataArray_44_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_12_MPORT_addr = replace_set;
  assign dataArray_44_12_MPORT_mask = _GEN_8592 & _GEN_7209;
  assign dataArray_44_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_13_cachedata_MPORT_en = dataArray_44_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_13_cachedata_MPORT_addr = dataArray_44_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_13_cachedata_MPORT_data = dataArray_44_13[dataArray_44_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_13_MPORT_addr = replace_set;
  assign dataArray_44_13_MPORT_mask = _GEN_8592 & _GEN_7211;
  assign dataArray_44_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_14_cachedata_MPORT_en = dataArray_44_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_14_cachedata_MPORT_addr = dataArray_44_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_14_cachedata_MPORT_data = dataArray_44_14[dataArray_44_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_14_MPORT_addr = replace_set;
  assign dataArray_44_14_MPORT_mask = _GEN_8592 & _GEN_7213;
  assign dataArray_44_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_44_15_cachedata_MPORT_en = dataArray_44_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_44_15_cachedata_MPORT_addr = dataArray_44_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_44_15_cachedata_MPORT_data = dataArray_44_15[dataArray_44_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_44_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_44_15_MPORT_addr = replace_set;
  assign dataArray_44_15_MPORT_mask = _GEN_8592 & _GEN_7215;
  assign dataArray_44_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_0_cachedata_MPORT_en = dataArray_45_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_0_cachedata_MPORT_addr = dataArray_45_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_0_cachedata_MPORT_data = dataArray_45_0[dataArray_45_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_0_MPORT_addr = replace_set;
  assign dataArray_45_0_MPORT_mask = _GEN_8624 & _GEN_7185;
  assign dataArray_45_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_1_cachedata_MPORT_en = dataArray_45_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_1_cachedata_MPORT_addr = dataArray_45_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_1_cachedata_MPORT_data = dataArray_45_1[dataArray_45_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_1_MPORT_addr = replace_set;
  assign dataArray_45_1_MPORT_mask = _GEN_8624 & _GEN_7187;
  assign dataArray_45_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_2_cachedata_MPORT_en = dataArray_45_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_2_cachedata_MPORT_addr = dataArray_45_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_2_cachedata_MPORT_data = dataArray_45_2[dataArray_45_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_2_MPORT_addr = replace_set;
  assign dataArray_45_2_MPORT_mask = _GEN_8624 & _GEN_7189;
  assign dataArray_45_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_3_cachedata_MPORT_en = dataArray_45_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_3_cachedata_MPORT_addr = dataArray_45_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_3_cachedata_MPORT_data = dataArray_45_3[dataArray_45_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_3_MPORT_addr = replace_set;
  assign dataArray_45_3_MPORT_mask = _GEN_8624 & _GEN_7191;
  assign dataArray_45_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_4_cachedata_MPORT_en = dataArray_45_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_4_cachedata_MPORT_addr = dataArray_45_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_4_cachedata_MPORT_data = dataArray_45_4[dataArray_45_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_4_MPORT_addr = replace_set;
  assign dataArray_45_4_MPORT_mask = _GEN_8624 & _GEN_7193;
  assign dataArray_45_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_5_cachedata_MPORT_en = dataArray_45_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_5_cachedata_MPORT_addr = dataArray_45_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_5_cachedata_MPORT_data = dataArray_45_5[dataArray_45_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_5_MPORT_addr = replace_set;
  assign dataArray_45_5_MPORT_mask = _GEN_8624 & _GEN_7195;
  assign dataArray_45_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_6_cachedata_MPORT_en = dataArray_45_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_6_cachedata_MPORT_addr = dataArray_45_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_6_cachedata_MPORT_data = dataArray_45_6[dataArray_45_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_6_MPORT_addr = replace_set;
  assign dataArray_45_6_MPORT_mask = _GEN_8624 & _GEN_7197;
  assign dataArray_45_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_7_cachedata_MPORT_en = dataArray_45_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_7_cachedata_MPORT_addr = dataArray_45_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_7_cachedata_MPORT_data = dataArray_45_7[dataArray_45_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_7_MPORT_addr = replace_set;
  assign dataArray_45_7_MPORT_mask = _GEN_8624 & _GEN_7199;
  assign dataArray_45_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_8_cachedata_MPORT_en = dataArray_45_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_8_cachedata_MPORT_addr = dataArray_45_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_8_cachedata_MPORT_data = dataArray_45_8[dataArray_45_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_8_MPORT_addr = replace_set;
  assign dataArray_45_8_MPORT_mask = _GEN_8624 & _GEN_7201;
  assign dataArray_45_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_9_cachedata_MPORT_en = dataArray_45_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_9_cachedata_MPORT_addr = dataArray_45_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_9_cachedata_MPORT_data = dataArray_45_9[dataArray_45_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_9_MPORT_addr = replace_set;
  assign dataArray_45_9_MPORT_mask = _GEN_8624 & _GEN_7203;
  assign dataArray_45_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_10_cachedata_MPORT_en = dataArray_45_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_10_cachedata_MPORT_addr = dataArray_45_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_10_cachedata_MPORT_data = dataArray_45_10[dataArray_45_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_10_MPORT_addr = replace_set;
  assign dataArray_45_10_MPORT_mask = _GEN_8624 & _GEN_7205;
  assign dataArray_45_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_11_cachedata_MPORT_en = dataArray_45_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_11_cachedata_MPORT_addr = dataArray_45_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_11_cachedata_MPORT_data = dataArray_45_11[dataArray_45_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_11_MPORT_addr = replace_set;
  assign dataArray_45_11_MPORT_mask = _GEN_8624 & _GEN_7207;
  assign dataArray_45_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_12_cachedata_MPORT_en = dataArray_45_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_12_cachedata_MPORT_addr = dataArray_45_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_12_cachedata_MPORT_data = dataArray_45_12[dataArray_45_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_12_MPORT_addr = replace_set;
  assign dataArray_45_12_MPORT_mask = _GEN_8624 & _GEN_7209;
  assign dataArray_45_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_13_cachedata_MPORT_en = dataArray_45_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_13_cachedata_MPORT_addr = dataArray_45_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_13_cachedata_MPORT_data = dataArray_45_13[dataArray_45_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_13_MPORT_addr = replace_set;
  assign dataArray_45_13_MPORT_mask = _GEN_8624 & _GEN_7211;
  assign dataArray_45_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_14_cachedata_MPORT_en = dataArray_45_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_14_cachedata_MPORT_addr = dataArray_45_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_14_cachedata_MPORT_data = dataArray_45_14[dataArray_45_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_14_MPORT_addr = replace_set;
  assign dataArray_45_14_MPORT_mask = _GEN_8624 & _GEN_7213;
  assign dataArray_45_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_45_15_cachedata_MPORT_en = dataArray_45_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_45_15_cachedata_MPORT_addr = dataArray_45_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_45_15_cachedata_MPORT_data = dataArray_45_15[dataArray_45_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_45_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_45_15_MPORT_addr = replace_set;
  assign dataArray_45_15_MPORT_mask = _GEN_8624 & _GEN_7215;
  assign dataArray_45_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_0_cachedata_MPORT_en = dataArray_46_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_0_cachedata_MPORT_addr = dataArray_46_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_0_cachedata_MPORT_data = dataArray_46_0[dataArray_46_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_0_MPORT_addr = replace_set;
  assign dataArray_46_0_MPORT_mask = _GEN_8656 & _GEN_7185;
  assign dataArray_46_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_1_cachedata_MPORT_en = dataArray_46_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_1_cachedata_MPORT_addr = dataArray_46_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_1_cachedata_MPORT_data = dataArray_46_1[dataArray_46_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_1_MPORT_addr = replace_set;
  assign dataArray_46_1_MPORT_mask = _GEN_8656 & _GEN_7187;
  assign dataArray_46_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_2_cachedata_MPORT_en = dataArray_46_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_2_cachedata_MPORT_addr = dataArray_46_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_2_cachedata_MPORT_data = dataArray_46_2[dataArray_46_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_2_MPORT_addr = replace_set;
  assign dataArray_46_2_MPORT_mask = _GEN_8656 & _GEN_7189;
  assign dataArray_46_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_3_cachedata_MPORT_en = dataArray_46_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_3_cachedata_MPORT_addr = dataArray_46_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_3_cachedata_MPORT_data = dataArray_46_3[dataArray_46_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_3_MPORT_addr = replace_set;
  assign dataArray_46_3_MPORT_mask = _GEN_8656 & _GEN_7191;
  assign dataArray_46_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_4_cachedata_MPORT_en = dataArray_46_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_4_cachedata_MPORT_addr = dataArray_46_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_4_cachedata_MPORT_data = dataArray_46_4[dataArray_46_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_4_MPORT_addr = replace_set;
  assign dataArray_46_4_MPORT_mask = _GEN_8656 & _GEN_7193;
  assign dataArray_46_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_5_cachedata_MPORT_en = dataArray_46_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_5_cachedata_MPORT_addr = dataArray_46_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_5_cachedata_MPORT_data = dataArray_46_5[dataArray_46_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_5_MPORT_addr = replace_set;
  assign dataArray_46_5_MPORT_mask = _GEN_8656 & _GEN_7195;
  assign dataArray_46_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_6_cachedata_MPORT_en = dataArray_46_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_6_cachedata_MPORT_addr = dataArray_46_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_6_cachedata_MPORT_data = dataArray_46_6[dataArray_46_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_6_MPORT_addr = replace_set;
  assign dataArray_46_6_MPORT_mask = _GEN_8656 & _GEN_7197;
  assign dataArray_46_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_7_cachedata_MPORT_en = dataArray_46_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_7_cachedata_MPORT_addr = dataArray_46_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_7_cachedata_MPORT_data = dataArray_46_7[dataArray_46_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_7_MPORT_addr = replace_set;
  assign dataArray_46_7_MPORT_mask = _GEN_8656 & _GEN_7199;
  assign dataArray_46_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_8_cachedata_MPORT_en = dataArray_46_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_8_cachedata_MPORT_addr = dataArray_46_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_8_cachedata_MPORT_data = dataArray_46_8[dataArray_46_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_8_MPORT_addr = replace_set;
  assign dataArray_46_8_MPORT_mask = _GEN_8656 & _GEN_7201;
  assign dataArray_46_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_9_cachedata_MPORT_en = dataArray_46_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_9_cachedata_MPORT_addr = dataArray_46_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_9_cachedata_MPORT_data = dataArray_46_9[dataArray_46_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_9_MPORT_addr = replace_set;
  assign dataArray_46_9_MPORT_mask = _GEN_8656 & _GEN_7203;
  assign dataArray_46_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_10_cachedata_MPORT_en = dataArray_46_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_10_cachedata_MPORT_addr = dataArray_46_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_10_cachedata_MPORT_data = dataArray_46_10[dataArray_46_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_10_MPORT_addr = replace_set;
  assign dataArray_46_10_MPORT_mask = _GEN_8656 & _GEN_7205;
  assign dataArray_46_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_11_cachedata_MPORT_en = dataArray_46_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_11_cachedata_MPORT_addr = dataArray_46_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_11_cachedata_MPORT_data = dataArray_46_11[dataArray_46_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_11_MPORT_addr = replace_set;
  assign dataArray_46_11_MPORT_mask = _GEN_8656 & _GEN_7207;
  assign dataArray_46_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_12_cachedata_MPORT_en = dataArray_46_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_12_cachedata_MPORT_addr = dataArray_46_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_12_cachedata_MPORT_data = dataArray_46_12[dataArray_46_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_12_MPORT_addr = replace_set;
  assign dataArray_46_12_MPORT_mask = _GEN_8656 & _GEN_7209;
  assign dataArray_46_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_13_cachedata_MPORT_en = dataArray_46_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_13_cachedata_MPORT_addr = dataArray_46_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_13_cachedata_MPORT_data = dataArray_46_13[dataArray_46_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_13_MPORT_addr = replace_set;
  assign dataArray_46_13_MPORT_mask = _GEN_8656 & _GEN_7211;
  assign dataArray_46_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_14_cachedata_MPORT_en = dataArray_46_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_14_cachedata_MPORT_addr = dataArray_46_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_14_cachedata_MPORT_data = dataArray_46_14[dataArray_46_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_14_MPORT_addr = replace_set;
  assign dataArray_46_14_MPORT_mask = _GEN_8656 & _GEN_7213;
  assign dataArray_46_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_46_15_cachedata_MPORT_en = dataArray_46_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_46_15_cachedata_MPORT_addr = dataArray_46_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_46_15_cachedata_MPORT_data = dataArray_46_15[dataArray_46_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_46_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_46_15_MPORT_addr = replace_set;
  assign dataArray_46_15_MPORT_mask = _GEN_8656 & _GEN_7215;
  assign dataArray_46_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_0_cachedata_MPORT_en = dataArray_47_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_0_cachedata_MPORT_addr = dataArray_47_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_0_cachedata_MPORT_data = dataArray_47_0[dataArray_47_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_0_MPORT_addr = replace_set;
  assign dataArray_47_0_MPORT_mask = _GEN_8688 & _GEN_7185;
  assign dataArray_47_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_1_cachedata_MPORT_en = dataArray_47_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_1_cachedata_MPORT_addr = dataArray_47_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_1_cachedata_MPORT_data = dataArray_47_1[dataArray_47_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_1_MPORT_addr = replace_set;
  assign dataArray_47_1_MPORT_mask = _GEN_8688 & _GEN_7187;
  assign dataArray_47_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_2_cachedata_MPORT_en = dataArray_47_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_2_cachedata_MPORT_addr = dataArray_47_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_2_cachedata_MPORT_data = dataArray_47_2[dataArray_47_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_2_MPORT_addr = replace_set;
  assign dataArray_47_2_MPORT_mask = _GEN_8688 & _GEN_7189;
  assign dataArray_47_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_3_cachedata_MPORT_en = dataArray_47_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_3_cachedata_MPORT_addr = dataArray_47_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_3_cachedata_MPORT_data = dataArray_47_3[dataArray_47_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_3_MPORT_addr = replace_set;
  assign dataArray_47_3_MPORT_mask = _GEN_8688 & _GEN_7191;
  assign dataArray_47_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_4_cachedata_MPORT_en = dataArray_47_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_4_cachedata_MPORT_addr = dataArray_47_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_4_cachedata_MPORT_data = dataArray_47_4[dataArray_47_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_4_MPORT_addr = replace_set;
  assign dataArray_47_4_MPORT_mask = _GEN_8688 & _GEN_7193;
  assign dataArray_47_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_5_cachedata_MPORT_en = dataArray_47_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_5_cachedata_MPORT_addr = dataArray_47_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_5_cachedata_MPORT_data = dataArray_47_5[dataArray_47_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_5_MPORT_addr = replace_set;
  assign dataArray_47_5_MPORT_mask = _GEN_8688 & _GEN_7195;
  assign dataArray_47_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_6_cachedata_MPORT_en = dataArray_47_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_6_cachedata_MPORT_addr = dataArray_47_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_6_cachedata_MPORT_data = dataArray_47_6[dataArray_47_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_6_MPORT_addr = replace_set;
  assign dataArray_47_6_MPORT_mask = _GEN_8688 & _GEN_7197;
  assign dataArray_47_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_7_cachedata_MPORT_en = dataArray_47_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_7_cachedata_MPORT_addr = dataArray_47_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_7_cachedata_MPORT_data = dataArray_47_7[dataArray_47_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_7_MPORT_addr = replace_set;
  assign dataArray_47_7_MPORT_mask = _GEN_8688 & _GEN_7199;
  assign dataArray_47_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_8_cachedata_MPORT_en = dataArray_47_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_8_cachedata_MPORT_addr = dataArray_47_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_8_cachedata_MPORT_data = dataArray_47_8[dataArray_47_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_8_MPORT_addr = replace_set;
  assign dataArray_47_8_MPORT_mask = _GEN_8688 & _GEN_7201;
  assign dataArray_47_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_9_cachedata_MPORT_en = dataArray_47_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_9_cachedata_MPORT_addr = dataArray_47_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_9_cachedata_MPORT_data = dataArray_47_9[dataArray_47_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_9_MPORT_addr = replace_set;
  assign dataArray_47_9_MPORT_mask = _GEN_8688 & _GEN_7203;
  assign dataArray_47_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_10_cachedata_MPORT_en = dataArray_47_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_10_cachedata_MPORT_addr = dataArray_47_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_10_cachedata_MPORT_data = dataArray_47_10[dataArray_47_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_10_MPORT_addr = replace_set;
  assign dataArray_47_10_MPORT_mask = _GEN_8688 & _GEN_7205;
  assign dataArray_47_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_11_cachedata_MPORT_en = dataArray_47_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_11_cachedata_MPORT_addr = dataArray_47_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_11_cachedata_MPORT_data = dataArray_47_11[dataArray_47_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_11_MPORT_addr = replace_set;
  assign dataArray_47_11_MPORT_mask = _GEN_8688 & _GEN_7207;
  assign dataArray_47_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_12_cachedata_MPORT_en = dataArray_47_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_12_cachedata_MPORT_addr = dataArray_47_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_12_cachedata_MPORT_data = dataArray_47_12[dataArray_47_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_12_MPORT_addr = replace_set;
  assign dataArray_47_12_MPORT_mask = _GEN_8688 & _GEN_7209;
  assign dataArray_47_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_13_cachedata_MPORT_en = dataArray_47_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_13_cachedata_MPORT_addr = dataArray_47_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_13_cachedata_MPORT_data = dataArray_47_13[dataArray_47_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_13_MPORT_addr = replace_set;
  assign dataArray_47_13_MPORT_mask = _GEN_8688 & _GEN_7211;
  assign dataArray_47_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_14_cachedata_MPORT_en = dataArray_47_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_14_cachedata_MPORT_addr = dataArray_47_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_14_cachedata_MPORT_data = dataArray_47_14[dataArray_47_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_14_MPORT_addr = replace_set;
  assign dataArray_47_14_MPORT_mask = _GEN_8688 & _GEN_7213;
  assign dataArray_47_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_47_15_cachedata_MPORT_en = dataArray_47_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_47_15_cachedata_MPORT_addr = dataArray_47_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_47_15_cachedata_MPORT_data = dataArray_47_15[dataArray_47_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_47_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_47_15_MPORT_addr = replace_set;
  assign dataArray_47_15_MPORT_mask = _GEN_8688 & _GEN_7215;
  assign dataArray_47_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_0_cachedata_MPORT_en = dataArray_48_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_0_cachedata_MPORT_addr = dataArray_48_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_0_cachedata_MPORT_data = dataArray_48_0[dataArray_48_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_0_MPORT_addr = replace_set;
  assign dataArray_48_0_MPORT_mask = _GEN_8720 & _GEN_7185;
  assign dataArray_48_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_1_cachedata_MPORT_en = dataArray_48_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_1_cachedata_MPORT_addr = dataArray_48_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_1_cachedata_MPORT_data = dataArray_48_1[dataArray_48_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_1_MPORT_addr = replace_set;
  assign dataArray_48_1_MPORT_mask = _GEN_8720 & _GEN_7187;
  assign dataArray_48_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_2_cachedata_MPORT_en = dataArray_48_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_2_cachedata_MPORT_addr = dataArray_48_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_2_cachedata_MPORT_data = dataArray_48_2[dataArray_48_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_2_MPORT_addr = replace_set;
  assign dataArray_48_2_MPORT_mask = _GEN_8720 & _GEN_7189;
  assign dataArray_48_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_3_cachedata_MPORT_en = dataArray_48_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_3_cachedata_MPORT_addr = dataArray_48_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_3_cachedata_MPORT_data = dataArray_48_3[dataArray_48_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_3_MPORT_addr = replace_set;
  assign dataArray_48_3_MPORT_mask = _GEN_8720 & _GEN_7191;
  assign dataArray_48_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_4_cachedata_MPORT_en = dataArray_48_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_4_cachedata_MPORT_addr = dataArray_48_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_4_cachedata_MPORT_data = dataArray_48_4[dataArray_48_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_4_MPORT_addr = replace_set;
  assign dataArray_48_4_MPORT_mask = _GEN_8720 & _GEN_7193;
  assign dataArray_48_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_5_cachedata_MPORT_en = dataArray_48_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_5_cachedata_MPORT_addr = dataArray_48_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_5_cachedata_MPORT_data = dataArray_48_5[dataArray_48_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_5_MPORT_addr = replace_set;
  assign dataArray_48_5_MPORT_mask = _GEN_8720 & _GEN_7195;
  assign dataArray_48_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_6_cachedata_MPORT_en = dataArray_48_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_6_cachedata_MPORT_addr = dataArray_48_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_6_cachedata_MPORT_data = dataArray_48_6[dataArray_48_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_6_MPORT_addr = replace_set;
  assign dataArray_48_6_MPORT_mask = _GEN_8720 & _GEN_7197;
  assign dataArray_48_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_7_cachedata_MPORT_en = dataArray_48_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_7_cachedata_MPORT_addr = dataArray_48_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_7_cachedata_MPORT_data = dataArray_48_7[dataArray_48_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_7_MPORT_addr = replace_set;
  assign dataArray_48_7_MPORT_mask = _GEN_8720 & _GEN_7199;
  assign dataArray_48_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_8_cachedata_MPORT_en = dataArray_48_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_8_cachedata_MPORT_addr = dataArray_48_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_8_cachedata_MPORT_data = dataArray_48_8[dataArray_48_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_8_MPORT_addr = replace_set;
  assign dataArray_48_8_MPORT_mask = _GEN_8720 & _GEN_7201;
  assign dataArray_48_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_9_cachedata_MPORT_en = dataArray_48_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_9_cachedata_MPORT_addr = dataArray_48_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_9_cachedata_MPORT_data = dataArray_48_9[dataArray_48_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_9_MPORT_addr = replace_set;
  assign dataArray_48_9_MPORT_mask = _GEN_8720 & _GEN_7203;
  assign dataArray_48_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_10_cachedata_MPORT_en = dataArray_48_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_10_cachedata_MPORT_addr = dataArray_48_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_10_cachedata_MPORT_data = dataArray_48_10[dataArray_48_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_10_MPORT_addr = replace_set;
  assign dataArray_48_10_MPORT_mask = _GEN_8720 & _GEN_7205;
  assign dataArray_48_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_11_cachedata_MPORT_en = dataArray_48_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_11_cachedata_MPORT_addr = dataArray_48_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_11_cachedata_MPORT_data = dataArray_48_11[dataArray_48_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_11_MPORT_addr = replace_set;
  assign dataArray_48_11_MPORT_mask = _GEN_8720 & _GEN_7207;
  assign dataArray_48_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_12_cachedata_MPORT_en = dataArray_48_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_12_cachedata_MPORT_addr = dataArray_48_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_12_cachedata_MPORT_data = dataArray_48_12[dataArray_48_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_12_MPORT_addr = replace_set;
  assign dataArray_48_12_MPORT_mask = _GEN_8720 & _GEN_7209;
  assign dataArray_48_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_13_cachedata_MPORT_en = dataArray_48_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_13_cachedata_MPORT_addr = dataArray_48_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_13_cachedata_MPORT_data = dataArray_48_13[dataArray_48_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_13_MPORT_addr = replace_set;
  assign dataArray_48_13_MPORT_mask = _GEN_8720 & _GEN_7211;
  assign dataArray_48_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_14_cachedata_MPORT_en = dataArray_48_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_14_cachedata_MPORT_addr = dataArray_48_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_14_cachedata_MPORT_data = dataArray_48_14[dataArray_48_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_14_MPORT_addr = replace_set;
  assign dataArray_48_14_MPORT_mask = _GEN_8720 & _GEN_7213;
  assign dataArray_48_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_48_15_cachedata_MPORT_en = dataArray_48_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_48_15_cachedata_MPORT_addr = dataArray_48_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_48_15_cachedata_MPORT_data = dataArray_48_15[dataArray_48_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_48_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_48_15_MPORT_addr = replace_set;
  assign dataArray_48_15_MPORT_mask = _GEN_8720 & _GEN_7215;
  assign dataArray_48_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_0_cachedata_MPORT_en = dataArray_49_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_0_cachedata_MPORT_addr = dataArray_49_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_0_cachedata_MPORT_data = dataArray_49_0[dataArray_49_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_0_MPORT_addr = replace_set;
  assign dataArray_49_0_MPORT_mask = _GEN_8752 & _GEN_7185;
  assign dataArray_49_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_1_cachedata_MPORT_en = dataArray_49_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_1_cachedata_MPORT_addr = dataArray_49_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_1_cachedata_MPORT_data = dataArray_49_1[dataArray_49_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_1_MPORT_addr = replace_set;
  assign dataArray_49_1_MPORT_mask = _GEN_8752 & _GEN_7187;
  assign dataArray_49_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_2_cachedata_MPORT_en = dataArray_49_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_2_cachedata_MPORT_addr = dataArray_49_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_2_cachedata_MPORT_data = dataArray_49_2[dataArray_49_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_2_MPORT_addr = replace_set;
  assign dataArray_49_2_MPORT_mask = _GEN_8752 & _GEN_7189;
  assign dataArray_49_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_3_cachedata_MPORT_en = dataArray_49_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_3_cachedata_MPORT_addr = dataArray_49_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_3_cachedata_MPORT_data = dataArray_49_3[dataArray_49_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_3_MPORT_addr = replace_set;
  assign dataArray_49_3_MPORT_mask = _GEN_8752 & _GEN_7191;
  assign dataArray_49_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_4_cachedata_MPORT_en = dataArray_49_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_4_cachedata_MPORT_addr = dataArray_49_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_4_cachedata_MPORT_data = dataArray_49_4[dataArray_49_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_4_MPORT_addr = replace_set;
  assign dataArray_49_4_MPORT_mask = _GEN_8752 & _GEN_7193;
  assign dataArray_49_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_5_cachedata_MPORT_en = dataArray_49_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_5_cachedata_MPORT_addr = dataArray_49_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_5_cachedata_MPORT_data = dataArray_49_5[dataArray_49_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_5_MPORT_addr = replace_set;
  assign dataArray_49_5_MPORT_mask = _GEN_8752 & _GEN_7195;
  assign dataArray_49_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_6_cachedata_MPORT_en = dataArray_49_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_6_cachedata_MPORT_addr = dataArray_49_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_6_cachedata_MPORT_data = dataArray_49_6[dataArray_49_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_6_MPORT_addr = replace_set;
  assign dataArray_49_6_MPORT_mask = _GEN_8752 & _GEN_7197;
  assign dataArray_49_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_7_cachedata_MPORT_en = dataArray_49_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_7_cachedata_MPORT_addr = dataArray_49_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_7_cachedata_MPORT_data = dataArray_49_7[dataArray_49_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_7_MPORT_addr = replace_set;
  assign dataArray_49_7_MPORT_mask = _GEN_8752 & _GEN_7199;
  assign dataArray_49_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_8_cachedata_MPORT_en = dataArray_49_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_8_cachedata_MPORT_addr = dataArray_49_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_8_cachedata_MPORT_data = dataArray_49_8[dataArray_49_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_8_MPORT_addr = replace_set;
  assign dataArray_49_8_MPORT_mask = _GEN_8752 & _GEN_7201;
  assign dataArray_49_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_9_cachedata_MPORT_en = dataArray_49_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_9_cachedata_MPORT_addr = dataArray_49_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_9_cachedata_MPORT_data = dataArray_49_9[dataArray_49_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_9_MPORT_addr = replace_set;
  assign dataArray_49_9_MPORT_mask = _GEN_8752 & _GEN_7203;
  assign dataArray_49_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_10_cachedata_MPORT_en = dataArray_49_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_10_cachedata_MPORT_addr = dataArray_49_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_10_cachedata_MPORT_data = dataArray_49_10[dataArray_49_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_10_MPORT_addr = replace_set;
  assign dataArray_49_10_MPORT_mask = _GEN_8752 & _GEN_7205;
  assign dataArray_49_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_11_cachedata_MPORT_en = dataArray_49_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_11_cachedata_MPORT_addr = dataArray_49_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_11_cachedata_MPORT_data = dataArray_49_11[dataArray_49_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_11_MPORT_addr = replace_set;
  assign dataArray_49_11_MPORT_mask = _GEN_8752 & _GEN_7207;
  assign dataArray_49_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_12_cachedata_MPORT_en = dataArray_49_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_12_cachedata_MPORT_addr = dataArray_49_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_12_cachedata_MPORT_data = dataArray_49_12[dataArray_49_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_12_MPORT_addr = replace_set;
  assign dataArray_49_12_MPORT_mask = _GEN_8752 & _GEN_7209;
  assign dataArray_49_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_13_cachedata_MPORT_en = dataArray_49_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_13_cachedata_MPORT_addr = dataArray_49_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_13_cachedata_MPORT_data = dataArray_49_13[dataArray_49_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_13_MPORT_addr = replace_set;
  assign dataArray_49_13_MPORT_mask = _GEN_8752 & _GEN_7211;
  assign dataArray_49_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_14_cachedata_MPORT_en = dataArray_49_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_14_cachedata_MPORT_addr = dataArray_49_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_14_cachedata_MPORT_data = dataArray_49_14[dataArray_49_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_14_MPORT_addr = replace_set;
  assign dataArray_49_14_MPORT_mask = _GEN_8752 & _GEN_7213;
  assign dataArray_49_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_49_15_cachedata_MPORT_en = dataArray_49_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_49_15_cachedata_MPORT_addr = dataArray_49_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_49_15_cachedata_MPORT_data = dataArray_49_15[dataArray_49_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_49_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_49_15_MPORT_addr = replace_set;
  assign dataArray_49_15_MPORT_mask = _GEN_8752 & _GEN_7215;
  assign dataArray_49_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_0_cachedata_MPORT_en = dataArray_50_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_0_cachedata_MPORT_addr = dataArray_50_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_0_cachedata_MPORT_data = dataArray_50_0[dataArray_50_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_0_MPORT_addr = replace_set;
  assign dataArray_50_0_MPORT_mask = _GEN_8784 & _GEN_7185;
  assign dataArray_50_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_1_cachedata_MPORT_en = dataArray_50_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_1_cachedata_MPORT_addr = dataArray_50_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_1_cachedata_MPORT_data = dataArray_50_1[dataArray_50_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_1_MPORT_addr = replace_set;
  assign dataArray_50_1_MPORT_mask = _GEN_8784 & _GEN_7187;
  assign dataArray_50_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_2_cachedata_MPORT_en = dataArray_50_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_2_cachedata_MPORT_addr = dataArray_50_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_2_cachedata_MPORT_data = dataArray_50_2[dataArray_50_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_2_MPORT_addr = replace_set;
  assign dataArray_50_2_MPORT_mask = _GEN_8784 & _GEN_7189;
  assign dataArray_50_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_3_cachedata_MPORT_en = dataArray_50_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_3_cachedata_MPORT_addr = dataArray_50_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_3_cachedata_MPORT_data = dataArray_50_3[dataArray_50_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_3_MPORT_addr = replace_set;
  assign dataArray_50_3_MPORT_mask = _GEN_8784 & _GEN_7191;
  assign dataArray_50_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_4_cachedata_MPORT_en = dataArray_50_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_4_cachedata_MPORT_addr = dataArray_50_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_4_cachedata_MPORT_data = dataArray_50_4[dataArray_50_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_4_MPORT_addr = replace_set;
  assign dataArray_50_4_MPORT_mask = _GEN_8784 & _GEN_7193;
  assign dataArray_50_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_5_cachedata_MPORT_en = dataArray_50_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_5_cachedata_MPORT_addr = dataArray_50_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_5_cachedata_MPORT_data = dataArray_50_5[dataArray_50_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_5_MPORT_addr = replace_set;
  assign dataArray_50_5_MPORT_mask = _GEN_8784 & _GEN_7195;
  assign dataArray_50_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_6_cachedata_MPORT_en = dataArray_50_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_6_cachedata_MPORT_addr = dataArray_50_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_6_cachedata_MPORT_data = dataArray_50_6[dataArray_50_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_6_MPORT_addr = replace_set;
  assign dataArray_50_6_MPORT_mask = _GEN_8784 & _GEN_7197;
  assign dataArray_50_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_7_cachedata_MPORT_en = dataArray_50_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_7_cachedata_MPORT_addr = dataArray_50_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_7_cachedata_MPORT_data = dataArray_50_7[dataArray_50_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_7_MPORT_addr = replace_set;
  assign dataArray_50_7_MPORT_mask = _GEN_8784 & _GEN_7199;
  assign dataArray_50_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_8_cachedata_MPORT_en = dataArray_50_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_8_cachedata_MPORT_addr = dataArray_50_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_8_cachedata_MPORT_data = dataArray_50_8[dataArray_50_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_8_MPORT_addr = replace_set;
  assign dataArray_50_8_MPORT_mask = _GEN_8784 & _GEN_7201;
  assign dataArray_50_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_9_cachedata_MPORT_en = dataArray_50_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_9_cachedata_MPORT_addr = dataArray_50_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_9_cachedata_MPORT_data = dataArray_50_9[dataArray_50_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_9_MPORT_addr = replace_set;
  assign dataArray_50_9_MPORT_mask = _GEN_8784 & _GEN_7203;
  assign dataArray_50_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_10_cachedata_MPORT_en = dataArray_50_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_10_cachedata_MPORT_addr = dataArray_50_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_10_cachedata_MPORT_data = dataArray_50_10[dataArray_50_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_10_MPORT_addr = replace_set;
  assign dataArray_50_10_MPORT_mask = _GEN_8784 & _GEN_7205;
  assign dataArray_50_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_11_cachedata_MPORT_en = dataArray_50_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_11_cachedata_MPORT_addr = dataArray_50_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_11_cachedata_MPORT_data = dataArray_50_11[dataArray_50_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_11_MPORT_addr = replace_set;
  assign dataArray_50_11_MPORT_mask = _GEN_8784 & _GEN_7207;
  assign dataArray_50_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_12_cachedata_MPORT_en = dataArray_50_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_12_cachedata_MPORT_addr = dataArray_50_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_12_cachedata_MPORT_data = dataArray_50_12[dataArray_50_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_12_MPORT_addr = replace_set;
  assign dataArray_50_12_MPORT_mask = _GEN_8784 & _GEN_7209;
  assign dataArray_50_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_13_cachedata_MPORT_en = dataArray_50_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_13_cachedata_MPORT_addr = dataArray_50_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_13_cachedata_MPORT_data = dataArray_50_13[dataArray_50_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_13_MPORT_addr = replace_set;
  assign dataArray_50_13_MPORT_mask = _GEN_8784 & _GEN_7211;
  assign dataArray_50_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_14_cachedata_MPORT_en = dataArray_50_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_14_cachedata_MPORT_addr = dataArray_50_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_14_cachedata_MPORT_data = dataArray_50_14[dataArray_50_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_14_MPORT_addr = replace_set;
  assign dataArray_50_14_MPORT_mask = _GEN_8784 & _GEN_7213;
  assign dataArray_50_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_50_15_cachedata_MPORT_en = dataArray_50_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_50_15_cachedata_MPORT_addr = dataArray_50_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_50_15_cachedata_MPORT_data = dataArray_50_15[dataArray_50_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_50_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_50_15_MPORT_addr = replace_set;
  assign dataArray_50_15_MPORT_mask = _GEN_8784 & _GEN_7215;
  assign dataArray_50_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_0_cachedata_MPORT_en = dataArray_51_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_0_cachedata_MPORT_addr = dataArray_51_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_0_cachedata_MPORT_data = dataArray_51_0[dataArray_51_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_0_MPORT_addr = replace_set;
  assign dataArray_51_0_MPORT_mask = _GEN_8816 & _GEN_7185;
  assign dataArray_51_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_1_cachedata_MPORT_en = dataArray_51_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_1_cachedata_MPORT_addr = dataArray_51_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_1_cachedata_MPORT_data = dataArray_51_1[dataArray_51_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_1_MPORT_addr = replace_set;
  assign dataArray_51_1_MPORT_mask = _GEN_8816 & _GEN_7187;
  assign dataArray_51_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_2_cachedata_MPORT_en = dataArray_51_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_2_cachedata_MPORT_addr = dataArray_51_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_2_cachedata_MPORT_data = dataArray_51_2[dataArray_51_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_2_MPORT_addr = replace_set;
  assign dataArray_51_2_MPORT_mask = _GEN_8816 & _GEN_7189;
  assign dataArray_51_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_3_cachedata_MPORT_en = dataArray_51_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_3_cachedata_MPORT_addr = dataArray_51_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_3_cachedata_MPORT_data = dataArray_51_3[dataArray_51_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_3_MPORT_addr = replace_set;
  assign dataArray_51_3_MPORT_mask = _GEN_8816 & _GEN_7191;
  assign dataArray_51_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_4_cachedata_MPORT_en = dataArray_51_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_4_cachedata_MPORT_addr = dataArray_51_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_4_cachedata_MPORT_data = dataArray_51_4[dataArray_51_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_4_MPORT_addr = replace_set;
  assign dataArray_51_4_MPORT_mask = _GEN_8816 & _GEN_7193;
  assign dataArray_51_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_5_cachedata_MPORT_en = dataArray_51_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_5_cachedata_MPORT_addr = dataArray_51_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_5_cachedata_MPORT_data = dataArray_51_5[dataArray_51_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_5_MPORT_addr = replace_set;
  assign dataArray_51_5_MPORT_mask = _GEN_8816 & _GEN_7195;
  assign dataArray_51_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_6_cachedata_MPORT_en = dataArray_51_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_6_cachedata_MPORT_addr = dataArray_51_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_6_cachedata_MPORT_data = dataArray_51_6[dataArray_51_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_6_MPORT_addr = replace_set;
  assign dataArray_51_6_MPORT_mask = _GEN_8816 & _GEN_7197;
  assign dataArray_51_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_7_cachedata_MPORT_en = dataArray_51_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_7_cachedata_MPORT_addr = dataArray_51_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_7_cachedata_MPORT_data = dataArray_51_7[dataArray_51_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_7_MPORT_addr = replace_set;
  assign dataArray_51_7_MPORT_mask = _GEN_8816 & _GEN_7199;
  assign dataArray_51_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_8_cachedata_MPORT_en = dataArray_51_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_8_cachedata_MPORT_addr = dataArray_51_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_8_cachedata_MPORT_data = dataArray_51_8[dataArray_51_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_8_MPORT_addr = replace_set;
  assign dataArray_51_8_MPORT_mask = _GEN_8816 & _GEN_7201;
  assign dataArray_51_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_9_cachedata_MPORT_en = dataArray_51_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_9_cachedata_MPORT_addr = dataArray_51_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_9_cachedata_MPORT_data = dataArray_51_9[dataArray_51_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_9_MPORT_addr = replace_set;
  assign dataArray_51_9_MPORT_mask = _GEN_8816 & _GEN_7203;
  assign dataArray_51_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_10_cachedata_MPORT_en = dataArray_51_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_10_cachedata_MPORT_addr = dataArray_51_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_10_cachedata_MPORT_data = dataArray_51_10[dataArray_51_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_10_MPORT_addr = replace_set;
  assign dataArray_51_10_MPORT_mask = _GEN_8816 & _GEN_7205;
  assign dataArray_51_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_11_cachedata_MPORT_en = dataArray_51_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_11_cachedata_MPORT_addr = dataArray_51_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_11_cachedata_MPORT_data = dataArray_51_11[dataArray_51_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_11_MPORT_addr = replace_set;
  assign dataArray_51_11_MPORT_mask = _GEN_8816 & _GEN_7207;
  assign dataArray_51_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_12_cachedata_MPORT_en = dataArray_51_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_12_cachedata_MPORT_addr = dataArray_51_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_12_cachedata_MPORT_data = dataArray_51_12[dataArray_51_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_12_MPORT_addr = replace_set;
  assign dataArray_51_12_MPORT_mask = _GEN_8816 & _GEN_7209;
  assign dataArray_51_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_13_cachedata_MPORT_en = dataArray_51_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_13_cachedata_MPORT_addr = dataArray_51_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_13_cachedata_MPORT_data = dataArray_51_13[dataArray_51_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_13_MPORT_addr = replace_set;
  assign dataArray_51_13_MPORT_mask = _GEN_8816 & _GEN_7211;
  assign dataArray_51_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_14_cachedata_MPORT_en = dataArray_51_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_14_cachedata_MPORT_addr = dataArray_51_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_14_cachedata_MPORT_data = dataArray_51_14[dataArray_51_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_14_MPORT_addr = replace_set;
  assign dataArray_51_14_MPORT_mask = _GEN_8816 & _GEN_7213;
  assign dataArray_51_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_51_15_cachedata_MPORT_en = dataArray_51_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_51_15_cachedata_MPORT_addr = dataArray_51_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_51_15_cachedata_MPORT_data = dataArray_51_15[dataArray_51_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_51_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_51_15_MPORT_addr = replace_set;
  assign dataArray_51_15_MPORT_mask = _GEN_8816 & _GEN_7215;
  assign dataArray_51_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_0_cachedata_MPORT_en = dataArray_52_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_0_cachedata_MPORT_addr = dataArray_52_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_0_cachedata_MPORT_data = dataArray_52_0[dataArray_52_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_0_MPORT_addr = replace_set;
  assign dataArray_52_0_MPORT_mask = _GEN_8848 & _GEN_7185;
  assign dataArray_52_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_1_cachedata_MPORT_en = dataArray_52_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_1_cachedata_MPORT_addr = dataArray_52_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_1_cachedata_MPORT_data = dataArray_52_1[dataArray_52_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_1_MPORT_addr = replace_set;
  assign dataArray_52_1_MPORT_mask = _GEN_8848 & _GEN_7187;
  assign dataArray_52_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_2_cachedata_MPORT_en = dataArray_52_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_2_cachedata_MPORT_addr = dataArray_52_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_2_cachedata_MPORT_data = dataArray_52_2[dataArray_52_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_2_MPORT_addr = replace_set;
  assign dataArray_52_2_MPORT_mask = _GEN_8848 & _GEN_7189;
  assign dataArray_52_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_3_cachedata_MPORT_en = dataArray_52_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_3_cachedata_MPORT_addr = dataArray_52_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_3_cachedata_MPORT_data = dataArray_52_3[dataArray_52_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_3_MPORT_addr = replace_set;
  assign dataArray_52_3_MPORT_mask = _GEN_8848 & _GEN_7191;
  assign dataArray_52_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_4_cachedata_MPORT_en = dataArray_52_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_4_cachedata_MPORT_addr = dataArray_52_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_4_cachedata_MPORT_data = dataArray_52_4[dataArray_52_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_4_MPORT_addr = replace_set;
  assign dataArray_52_4_MPORT_mask = _GEN_8848 & _GEN_7193;
  assign dataArray_52_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_5_cachedata_MPORT_en = dataArray_52_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_5_cachedata_MPORT_addr = dataArray_52_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_5_cachedata_MPORT_data = dataArray_52_5[dataArray_52_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_5_MPORT_addr = replace_set;
  assign dataArray_52_5_MPORT_mask = _GEN_8848 & _GEN_7195;
  assign dataArray_52_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_6_cachedata_MPORT_en = dataArray_52_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_6_cachedata_MPORT_addr = dataArray_52_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_6_cachedata_MPORT_data = dataArray_52_6[dataArray_52_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_6_MPORT_addr = replace_set;
  assign dataArray_52_6_MPORT_mask = _GEN_8848 & _GEN_7197;
  assign dataArray_52_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_7_cachedata_MPORT_en = dataArray_52_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_7_cachedata_MPORT_addr = dataArray_52_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_7_cachedata_MPORT_data = dataArray_52_7[dataArray_52_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_7_MPORT_addr = replace_set;
  assign dataArray_52_7_MPORT_mask = _GEN_8848 & _GEN_7199;
  assign dataArray_52_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_8_cachedata_MPORT_en = dataArray_52_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_8_cachedata_MPORT_addr = dataArray_52_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_8_cachedata_MPORT_data = dataArray_52_8[dataArray_52_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_8_MPORT_addr = replace_set;
  assign dataArray_52_8_MPORT_mask = _GEN_8848 & _GEN_7201;
  assign dataArray_52_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_9_cachedata_MPORT_en = dataArray_52_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_9_cachedata_MPORT_addr = dataArray_52_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_9_cachedata_MPORT_data = dataArray_52_9[dataArray_52_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_9_MPORT_addr = replace_set;
  assign dataArray_52_9_MPORT_mask = _GEN_8848 & _GEN_7203;
  assign dataArray_52_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_10_cachedata_MPORT_en = dataArray_52_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_10_cachedata_MPORT_addr = dataArray_52_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_10_cachedata_MPORT_data = dataArray_52_10[dataArray_52_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_10_MPORT_addr = replace_set;
  assign dataArray_52_10_MPORT_mask = _GEN_8848 & _GEN_7205;
  assign dataArray_52_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_11_cachedata_MPORT_en = dataArray_52_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_11_cachedata_MPORT_addr = dataArray_52_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_11_cachedata_MPORT_data = dataArray_52_11[dataArray_52_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_11_MPORT_addr = replace_set;
  assign dataArray_52_11_MPORT_mask = _GEN_8848 & _GEN_7207;
  assign dataArray_52_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_12_cachedata_MPORT_en = dataArray_52_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_12_cachedata_MPORT_addr = dataArray_52_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_12_cachedata_MPORT_data = dataArray_52_12[dataArray_52_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_12_MPORT_addr = replace_set;
  assign dataArray_52_12_MPORT_mask = _GEN_8848 & _GEN_7209;
  assign dataArray_52_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_13_cachedata_MPORT_en = dataArray_52_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_13_cachedata_MPORT_addr = dataArray_52_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_13_cachedata_MPORT_data = dataArray_52_13[dataArray_52_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_13_MPORT_addr = replace_set;
  assign dataArray_52_13_MPORT_mask = _GEN_8848 & _GEN_7211;
  assign dataArray_52_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_14_cachedata_MPORT_en = dataArray_52_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_14_cachedata_MPORT_addr = dataArray_52_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_14_cachedata_MPORT_data = dataArray_52_14[dataArray_52_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_14_MPORT_addr = replace_set;
  assign dataArray_52_14_MPORT_mask = _GEN_8848 & _GEN_7213;
  assign dataArray_52_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_52_15_cachedata_MPORT_en = dataArray_52_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_52_15_cachedata_MPORT_addr = dataArray_52_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_52_15_cachedata_MPORT_data = dataArray_52_15[dataArray_52_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_52_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_52_15_MPORT_addr = replace_set;
  assign dataArray_52_15_MPORT_mask = _GEN_8848 & _GEN_7215;
  assign dataArray_52_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_0_cachedata_MPORT_en = dataArray_53_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_0_cachedata_MPORT_addr = dataArray_53_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_0_cachedata_MPORT_data = dataArray_53_0[dataArray_53_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_0_MPORT_addr = replace_set;
  assign dataArray_53_0_MPORT_mask = _GEN_8880 & _GEN_7185;
  assign dataArray_53_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_1_cachedata_MPORT_en = dataArray_53_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_1_cachedata_MPORT_addr = dataArray_53_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_1_cachedata_MPORT_data = dataArray_53_1[dataArray_53_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_1_MPORT_addr = replace_set;
  assign dataArray_53_1_MPORT_mask = _GEN_8880 & _GEN_7187;
  assign dataArray_53_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_2_cachedata_MPORT_en = dataArray_53_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_2_cachedata_MPORT_addr = dataArray_53_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_2_cachedata_MPORT_data = dataArray_53_2[dataArray_53_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_2_MPORT_addr = replace_set;
  assign dataArray_53_2_MPORT_mask = _GEN_8880 & _GEN_7189;
  assign dataArray_53_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_3_cachedata_MPORT_en = dataArray_53_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_3_cachedata_MPORT_addr = dataArray_53_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_3_cachedata_MPORT_data = dataArray_53_3[dataArray_53_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_3_MPORT_addr = replace_set;
  assign dataArray_53_3_MPORT_mask = _GEN_8880 & _GEN_7191;
  assign dataArray_53_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_4_cachedata_MPORT_en = dataArray_53_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_4_cachedata_MPORT_addr = dataArray_53_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_4_cachedata_MPORT_data = dataArray_53_4[dataArray_53_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_4_MPORT_addr = replace_set;
  assign dataArray_53_4_MPORT_mask = _GEN_8880 & _GEN_7193;
  assign dataArray_53_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_5_cachedata_MPORT_en = dataArray_53_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_5_cachedata_MPORT_addr = dataArray_53_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_5_cachedata_MPORT_data = dataArray_53_5[dataArray_53_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_5_MPORT_addr = replace_set;
  assign dataArray_53_5_MPORT_mask = _GEN_8880 & _GEN_7195;
  assign dataArray_53_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_6_cachedata_MPORT_en = dataArray_53_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_6_cachedata_MPORT_addr = dataArray_53_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_6_cachedata_MPORT_data = dataArray_53_6[dataArray_53_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_6_MPORT_addr = replace_set;
  assign dataArray_53_6_MPORT_mask = _GEN_8880 & _GEN_7197;
  assign dataArray_53_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_7_cachedata_MPORT_en = dataArray_53_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_7_cachedata_MPORT_addr = dataArray_53_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_7_cachedata_MPORT_data = dataArray_53_7[dataArray_53_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_7_MPORT_addr = replace_set;
  assign dataArray_53_7_MPORT_mask = _GEN_8880 & _GEN_7199;
  assign dataArray_53_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_8_cachedata_MPORT_en = dataArray_53_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_8_cachedata_MPORT_addr = dataArray_53_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_8_cachedata_MPORT_data = dataArray_53_8[dataArray_53_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_8_MPORT_addr = replace_set;
  assign dataArray_53_8_MPORT_mask = _GEN_8880 & _GEN_7201;
  assign dataArray_53_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_9_cachedata_MPORT_en = dataArray_53_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_9_cachedata_MPORT_addr = dataArray_53_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_9_cachedata_MPORT_data = dataArray_53_9[dataArray_53_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_9_MPORT_addr = replace_set;
  assign dataArray_53_9_MPORT_mask = _GEN_8880 & _GEN_7203;
  assign dataArray_53_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_10_cachedata_MPORT_en = dataArray_53_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_10_cachedata_MPORT_addr = dataArray_53_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_10_cachedata_MPORT_data = dataArray_53_10[dataArray_53_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_10_MPORT_addr = replace_set;
  assign dataArray_53_10_MPORT_mask = _GEN_8880 & _GEN_7205;
  assign dataArray_53_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_11_cachedata_MPORT_en = dataArray_53_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_11_cachedata_MPORT_addr = dataArray_53_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_11_cachedata_MPORT_data = dataArray_53_11[dataArray_53_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_11_MPORT_addr = replace_set;
  assign dataArray_53_11_MPORT_mask = _GEN_8880 & _GEN_7207;
  assign dataArray_53_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_12_cachedata_MPORT_en = dataArray_53_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_12_cachedata_MPORT_addr = dataArray_53_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_12_cachedata_MPORT_data = dataArray_53_12[dataArray_53_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_12_MPORT_addr = replace_set;
  assign dataArray_53_12_MPORT_mask = _GEN_8880 & _GEN_7209;
  assign dataArray_53_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_13_cachedata_MPORT_en = dataArray_53_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_13_cachedata_MPORT_addr = dataArray_53_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_13_cachedata_MPORT_data = dataArray_53_13[dataArray_53_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_13_MPORT_addr = replace_set;
  assign dataArray_53_13_MPORT_mask = _GEN_8880 & _GEN_7211;
  assign dataArray_53_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_14_cachedata_MPORT_en = dataArray_53_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_14_cachedata_MPORT_addr = dataArray_53_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_14_cachedata_MPORT_data = dataArray_53_14[dataArray_53_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_14_MPORT_addr = replace_set;
  assign dataArray_53_14_MPORT_mask = _GEN_8880 & _GEN_7213;
  assign dataArray_53_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_53_15_cachedata_MPORT_en = dataArray_53_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_53_15_cachedata_MPORT_addr = dataArray_53_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_53_15_cachedata_MPORT_data = dataArray_53_15[dataArray_53_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_53_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_53_15_MPORT_addr = replace_set;
  assign dataArray_53_15_MPORT_mask = _GEN_8880 & _GEN_7215;
  assign dataArray_53_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_0_cachedata_MPORT_en = dataArray_54_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_0_cachedata_MPORT_addr = dataArray_54_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_0_cachedata_MPORT_data = dataArray_54_0[dataArray_54_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_0_MPORT_addr = replace_set;
  assign dataArray_54_0_MPORT_mask = _GEN_8912 & _GEN_7185;
  assign dataArray_54_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_1_cachedata_MPORT_en = dataArray_54_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_1_cachedata_MPORT_addr = dataArray_54_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_1_cachedata_MPORT_data = dataArray_54_1[dataArray_54_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_1_MPORT_addr = replace_set;
  assign dataArray_54_1_MPORT_mask = _GEN_8912 & _GEN_7187;
  assign dataArray_54_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_2_cachedata_MPORT_en = dataArray_54_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_2_cachedata_MPORT_addr = dataArray_54_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_2_cachedata_MPORT_data = dataArray_54_2[dataArray_54_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_2_MPORT_addr = replace_set;
  assign dataArray_54_2_MPORT_mask = _GEN_8912 & _GEN_7189;
  assign dataArray_54_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_3_cachedata_MPORT_en = dataArray_54_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_3_cachedata_MPORT_addr = dataArray_54_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_3_cachedata_MPORT_data = dataArray_54_3[dataArray_54_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_3_MPORT_addr = replace_set;
  assign dataArray_54_3_MPORT_mask = _GEN_8912 & _GEN_7191;
  assign dataArray_54_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_4_cachedata_MPORT_en = dataArray_54_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_4_cachedata_MPORT_addr = dataArray_54_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_4_cachedata_MPORT_data = dataArray_54_4[dataArray_54_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_4_MPORT_addr = replace_set;
  assign dataArray_54_4_MPORT_mask = _GEN_8912 & _GEN_7193;
  assign dataArray_54_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_5_cachedata_MPORT_en = dataArray_54_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_5_cachedata_MPORT_addr = dataArray_54_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_5_cachedata_MPORT_data = dataArray_54_5[dataArray_54_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_5_MPORT_addr = replace_set;
  assign dataArray_54_5_MPORT_mask = _GEN_8912 & _GEN_7195;
  assign dataArray_54_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_6_cachedata_MPORT_en = dataArray_54_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_6_cachedata_MPORT_addr = dataArray_54_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_6_cachedata_MPORT_data = dataArray_54_6[dataArray_54_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_6_MPORT_addr = replace_set;
  assign dataArray_54_6_MPORT_mask = _GEN_8912 & _GEN_7197;
  assign dataArray_54_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_7_cachedata_MPORT_en = dataArray_54_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_7_cachedata_MPORT_addr = dataArray_54_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_7_cachedata_MPORT_data = dataArray_54_7[dataArray_54_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_7_MPORT_addr = replace_set;
  assign dataArray_54_7_MPORT_mask = _GEN_8912 & _GEN_7199;
  assign dataArray_54_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_8_cachedata_MPORT_en = dataArray_54_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_8_cachedata_MPORT_addr = dataArray_54_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_8_cachedata_MPORT_data = dataArray_54_8[dataArray_54_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_8_MPORT_addr = replace_set;
  assign dataArray_54_8_MPORT_mask = _GEN_8912 & _GEN_7201;
  assign dataArray_54_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_9_cachedata_MPORT_en = dataArray_54_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_9_cachedata_MPORT_addr = dataArray_54_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_9_cachedata_MPORT_data = dataArray_54_9[dataArray_54_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_9_MPORT_addr = replace_set;
  assign dataArray_54_9_MPORT_mask = _GEN_8912 & _GEN_7203;
  assign dataArray_54_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_10_cachedata_MPORT_en = dataArray_54_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_10_cachedata_MPORT_addr = dataArray_54_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_10_cachedata_MPORT_data = dataArray_54_10[dataArray_54_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_10_MPORT_addr = replace_set;
  assign dataArray_54_10_MPORT_mask = _GEN_8912 & _GEN_7205;
  assign dataArray_54_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_11_cachedata_MPORT_en = dataArray_54_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_11_cachedata_MPORT_addr = dataArray_54_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_11_cachedata_MPORT_data = dataArray_54_11[dataArray_54_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_11_MPORT_addr = replace_set;
  assign dataArray_54_11_MPORT_mask = _GEN_8912 & _GEN_7207;
  assign dataArray_54_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_12_cachedata_MPORT_en = dataArray_54_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_12_cachedata_MPORT_addr = dataArray_54_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_12_cachedata_MPORT_data = dataArray_54_12[dataArray_54_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_12_MPORT_addr = replace_set;
  assign dataArray_54_12_MPORT_mask = _GEN_8912 & _GEN_7209;
  assign dataArray_54_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_13_cachedata_MPORT_en = dataArray_54_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_13_cachedata_MPORT_addr = dataArray_54_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_13_cachedata_MPORT_data = dataArray_54_13[dataArray_54_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_13_MPORT_addr = replace_set;
  assign dataArray_54_13_MPORT_mask = _GEN_8912 & _GEN_7211;
  assign dataArray_54_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_14_cachedata_MPORT_en = dataArray_54_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_14_cachedata_MPORT_addr = dataArray_54_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_14_cachedata_MPORT_data = dataArray_54_14[dataArray_54_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_14_MPORT_addr = replace_set;
  assign dataArray_54_14_MPORT_mask = _GEN_8912 & _GEN_7213;
  assign dataArray_54_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_54_15_cachedata_MPORT_en = dataArray_54_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_54_15_cachedata_MPORT_addr = dataArray_54_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_54_15_cachedata_MPORT_data = dataArray_54_15[dataArray_54_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_54_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_54_15_MPORT_addr = replace_set;
  assign dataArray_54_15_MPORT_mask = _GEN_8912 & _GEN_7215;
  assign dataArray_54_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_0_cachedata_MPORT_en = dataArray_55_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_0_cachedata_MPORT_addr = dataArray_55_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_0_cachedata_MPORT_data = dataArray_55_0[dataArray_55_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_0_MPORT_addr = replace_set;
  assign dataArray_55_0_MPORT_mask = _GEN_8944 & _GEN_7185;
  assign dataArray_55_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_1_cachedata_MPORT_en = dataArray_55_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_1_cachedata_MPORT_addr = dataArray_55_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_1_cachedata_MPORT_data = dataArray_55_1[dataArray_55_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_1_MPORT_addr = replace_set;
  assign dataArray_55_1_MPORT_mask = _GEN_8944 & _GEN_7187;
  assign dataArray_55_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_2_cachedata_MPORT_en = dataArray_55_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_2_cachedata_MPORT_addr = dataArray_55_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_2_cachedata_MPORT_data = dataArray_55_2[dataArray_55_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_2_MPORT_addr = replace_set;
  assign dataArray_55_2_MPORT_mask = _GEN_8944 & _GEN_7189;
  assign dataArray_55_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_3_cachedata_MPORT_en = dataArray_55_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_3_cachedata_MPORT_addr = dataArray_55_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_3_cachedata_MPORT_data = dataArray_55_3[dataArray_55_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_3_MPORT_addr = replace_set;
  assign dataArray_55_3_MPORT_mask = _GEN_8944 & _GEN_7191;
  assign dataArray_55_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_4_cachedata_MPORT_en = dataArray_55_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_4_cachedata_MPORT_addr = dataArray_55_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_4_cachedata_MPORT_data = dataArray_55_4[dataArray_55_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_4_MPORT_addr = replace_set;
  assign dataArray_55_4_MPORT_mask = _GEN_8944 & _GEN_7193;
  assign dataArray_55_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_5_cachedata_MPORT_en = dataArray_55_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_5_cachedata_MPORT_addr = dataArray_55_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_5_cachedata_MPORT_data = dataArray_55_5[dataArray_55_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_5_MPORT_addr = replace_set;
  assign dataArray_55_5_MPORT_mask = _GEN_8944 & _GEN_7195;
  assign dataArray_55_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_6_cachedata_MPORT_en = dataArray_55_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_6_cachedata_MPORT_addr = dataArray_55_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_6_cachedata_MPORT_data = dataArray_55_6[dataArray_55_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_6_MPORT_addr = replace_set;
  assign dataArray_55_6_MPORT_mask = _GEN_8944 & _GEN_7197;
  assign dataArray_55_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_7_cachedata_MPORT_en = dataArray_55_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_7_cachedata_MPORT_addr = dataArray_55_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_7_cachedata_MPORT_data = dataArray_55_7[dataArray_55_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_7_MPORT_addr = replace_set;
  assign dataArray_55_7_MPORT_mask = _GEN_8944 & _GEN_7199;
  assign dataArray_55_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_8_cachedata_MPORT_en = dataArray_55_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_8_cachedata_MPORT_addr = dataArray_55_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_8_cachedata_MPORT_data = dataArray_55_8[dataArray_55_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_8_MPORT_addr = replace_set;
  assign dataArray_55_8_MPORT_mask = _GEN_8944 & _GEN_7201;
  assign dataArray_55_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_9_cachedata_MPORT_en = dataArray_55_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_9_cachedata_MPORT_addr = dataArray_55_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_9_cachedata_MPORT_data = dataArray_55_9[dataArray_55_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_9_MPORT_addr = replace_set;
  assign dataArray_55_9_MPORT_mask = _GEN_8944 & _GEN_7203;
  assign dataArray_55_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_10_cachedata_MPORT_en = dataArray_55_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_10_cachedata_MPORT_addr = dataArray_55_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_10_cachedata_MPORT_data = dataArray_55_10[dataArray_55_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_10_MPORT_addr = replace_set;
  assign dataArray_55_10_MPORT_mask = _GEN_8944 & _GEN_7205;
  assign dataArray_55_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_11_cachedata_MPORT_en = dataArray_55_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_11_cachedata_MPORT_addr = dataArray_55_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_11_cachedata_MPORT_data = dataArray_55_11[dataArray_55_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_11_MPORT_addr = replace_set;
  assign dataArray_55_11_MPORT_mask = _GEN_8944 & _GEN_7207;
  assign dataArray_55_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_12_cachedata_MPORT_en = dataArray_55_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_12_cachedata_MPORT_addr = dataArray_55_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_12_cachedata_MPORT_data = dataArray_55_12[dataArray_55_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_12_MPORT_addr = replace_set;
  assign dataArray_55_12_MPORT_mask = _GEN_8944 & _GEN_7209;
  assign dataArray_55_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_13_cachedata_MPORT_en = dataArray_55_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_13_cachedata_MPORT_addr = dataArray_55_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_13_cachedata_MPORT_data = dataArray_55_13[dataArray_55_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_13_MPORT_addr = replace_set;
  assign dataArray_55_13_MPORT_mask = _GEN_8944 & _GEN_7211;
  assign dataArray_55_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_14_cachedata_MPORT_en = dataArray_55_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_14_cachedata_MPORT_addr = dataArray_55_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_14_cachedata_MPORT_data = dataArray_55_14[dataArray_55_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_14_MPORT_addr = replace_set;
  assign dataArray_55_14_MPORT_mask = _GEN_8944 & _GEN_7213;
  assign dataArray_55_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_55_15_cachedata_MPORT_en = dataArray_55_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_55_15_cachedata_MPORT_addr = dataArray_55_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_55_15_cachedata_MPORT_data = dataArray_55_15[dataArray_55_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_55_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_55_15_MPORT_addr = replace_set;
  assign dataArray_55_15_MPORT_mask = _GEN_8944 & _GEN_7215;
  assign dataArray_55_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_0_cachedata_MPORT_en = dataArray_56_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_0_cachedata_MPORT_addr = dataArray_56_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_0_cachedata_MPORT_data = dataArray_56_0[dataArray_56_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_0_MPORT_addr = replace_set;
  assign dataArray_56_0_MPORT_mask = _GEN_8976 & _GEN_7185;
  assign dataArray_56_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_1_cachedata_MPORT_en = dataArray_56_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_1_cachedata_MPORT_addr = dataArray_56_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_1_cachedata_MPORT_data = dataArray_56_1[dataArray_56_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_1_MPORT_addr = replace_set;
  assign dataArray_56_1_MPORT_mask = _GEN_8976 & _GEN_7187;
  assign dataArray_56_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_2_cachedata_MPORT_en = dataArray_56_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_2_cachedata_MPORT_addr = dataArray_56_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_2_cachedata_MPORT_data = dataArray_56_2[dataArray_56_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_2_MPORT_addr = replace_set;
  assign dataArray_56_2_MPORT_mask = _GEN_8976 & _GEN_7189;
  assign dataArray_56_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_3_cachedata_MPORT_en = dataArray_56_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_3_cachedata_MPORT_addr = dataArray_56_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_3_cachedata_MPORT_data = dataArray_56_3[dataArray_56_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_3_MPORT_addr = replace_set;
  assign dataArray_56_3_MPORT_mask = _GEN_8976 & _GEN_7191;
  assign dataArray_56_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_4_cachedata_MPORT_en = dataArray_56_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_4_cachedata_MPORT_addr = dataArray_56_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_4_cachedata_MPORT_data = dataArray_56_4[dataArray_56_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_4_MPORT_addr = replace_set;
  assign dataArray_56_4_MPORT_mask = _GEN_8976 & _GEN_7193;
  assign dataArray_56_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_5_cachedata_MPORT_en = dataArray_56_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_5_cachedata_MPORT_addr = dataArray_56_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_5_cachedata_MPORT_data = dataArray_56_5[dataArray_56_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_5_MPORT_addr = replace_set;
  assign dataArray_56_5_MPORT_mask = _GEN_8976 & _GEN_7195;
  assign dataArray_56_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_6_cachedata_MPORT_en = dataArray_56_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_6_cachedata_MPORT_addr = dataArray_56_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_6_cachedata_MPORT_data = dataArray_56_6[dataArray_56_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_6_MPORT_addr = replace_set;
  assign dataArray_56_6_MPORT_mask = _GEN_8976 & _GEN_7197;
  assign dataArray_56_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_7_cachedata_MPORT_en = dataArray_56_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_7_cachedata_MPORT_addr = dataArray_56_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_7_cachedata_MPORT_data = dataArray_56_7[dataArray_56_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_7_MPORT_addr = replace_set;
  assign dataArray_56_7_MPORT_mask = _GEN_8976 & _GEN_7199;
  assign dataArray_56_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_8_cachedata_MPORT_en = dataArray_56_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_8_cachedata_MPORT_addr = dataArray_56_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_8_cachedata_MPORT_data = dataArray_56_8[dataArray_56_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_8_MPORT_addr = replace_set;
  assign dataArray_56_8_MPORT_mask = _GEN_8976 & _GEN_7201;
  assign dataArray_56_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_9_cachedata_MPORT_en = dataArray_56_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_9_cachedata_MPORT_addr = dataArray_56_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_9_cachedata_MPORT_data = dataArray_56_9[dataArray_56_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_9_MPORT_addr = replace_set;
  assign dataArray_56_9_MPORT_mask = _GEN_8976 & _GEN_7203;
  assign dataArray_56_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_10_cachedata_MPORT_en = dataArray_56_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_10_cachedata_MPORT_addr = dataArray_56_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_10_cachedata_MPORT_data = dataArray_56_10[dataArray_56_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_10_MPORT_addr = replace_set;
  assign dataArray_56_10_MPORT_mask = _GEN_8976 & _GEN_7205;
  assign dataArray_56_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_11_cachedata_MPORT_en = dataArray_56_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_11_cachedata_MPORT_addr = dataArray_56_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_11_cachedata_MPORT_data = dataArray_56_11[dataArray_56_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_11_MPORT_addr = replace_set;
  assign dataArray_56_11_MPORT_mask = _GEN_8976 & _GEN_7207;
  assign dataArray_56_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_12_cachedata_MPORT_en = dataArray_56_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_12_cachedata_MPORT_addr = dataArray_56_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_12_cachedata_MPORT_data = dataArray_56_12[dataArray_56_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_12_MPORT_addr = replace_set;
  assign dataArray_56_12_MPORT_mask = _GEN_8976 & _GEN_7209;
  assign dataArray_56_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_13_cachedata_MPORT_en = dataArray_56_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_13_cachedata_MPORT_addr = dataArray_56_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_13_cachedata_MPORT_data = dataArray_56_13[dataArray_56_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_13_MPORT_addr = replace_set;
  assign dataArray_56_13_MPORT_mask = _GEN_8976 & _GEN_7211;
  assign dataArray_56_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_14_cachedata_MPORT_en = dataArray_56_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_14_cachedata_MPORT_addr = dataArray_56_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_14_cachedata_MPORT_data = dataArray_56_14[dataArray_56_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_14_MPORT_addr = replace_set;
  assign dataArray_56_14_MPORT_mask = _GEN_8976 & _GEN_7213;
  assign dataArray_56_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_56_15_cachedata_MPORT_en = dataArray_56_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_56_15_cachedata_MPORT_addr = dataArray_56_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_56_15_cachedata_MPORT_data = dataArray_56_15[dataArray_56_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_56_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_56_15_MPORT_addr = replace_set;
  assign dataArray_56_15_MPORT_mask = _GEN_8976 & _GEN_7215;
  assign dataArray_56_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_0_cachedata_MPORT_en = dataArray_57_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_0_cachedata_MPORT_addr = dataArray_57_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_0_cachedata_MPORT_data = dataArray_57_0[dataArray_57_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_0_MPORT_addr = replace_set;
  assign dataArray_57_0_MPORT_mask = _GEN_9008 & _GEN_7185;
  assign dataArray_57_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_1_cachedata_MPORT_en = dataArray_57_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_1_cachedata_MPORT_addr = dataArray_57_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_1_cachedata_MPORT_data = dataArray_57_1[dataArray_57_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_1_MPORT_addr = replace_set;
  assign dataArray_57_1_MPORT_mask = _GEN_9008 & _GEN_7187;
  assign dataArray_57_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_2_cachedata_MPORT_en = dataArray_57_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_2_cachedata_MPORT_addr = dataArray_57_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_2_cachedata_MPORT_data = dataArray_57_2[dataArray_57_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_2_MPORT_addr = replace_set;
  assign dataArray_57_2_MPORT_mask = _GEN_9008 & _GEN_7189;
  assign dataArray_57_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_3_cachedata_MPORT_en = dataArray_57_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_3_cachedata_MPORT_addr = dataArray_57_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_3_cachedata_MPORT_data = dataArray_57_3[dataArray_57_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_3_MPORT_addr = replace_set;
  assign dataArray_57_3_MPORT_mask = _GEN_9008 & _GEN_7191;
  assign dataArray_57_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_4_cachedata_MPORT_en = dataArray_57_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_4_cachedata_MPORT_addr = dataArray_57_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_4_cachedata_MPORT_data = dataArray_57_4[dataArray_57_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_4_MPORT_addr = replace_set;
  assign dataArray_57_4_MPORT_mask = _GEN_9008 & _GEN_7193;
  assign dataArray_57_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_5_cachedata_MPORT_en = dataArray_57_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_5_cachedata_MPORT_addr = dataArray_57_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_5_cachedata_MPORT_data = dataArray_57_5[dataArray_57_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_5_MPORT_addr = replace_set;
  assign dataArray_57_5_MPORT_mask = _GEN_9008 & _GEN_7195;
  assign dataArray_57_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_6_cachedata_MPORT_en = dataArray_57_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_6_cachedata_MPORT_addr = dataArray_57_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_6_cachedata_MPORT_data = dataArray_57_6[dataArray_57_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_6_MPORT_addr = replace_set;
  assign dataArray_57_6_MPORT_mask = _GEN_9008 & _GEN_7197;
  assign dataArray_57_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_7_cachedata_MPORT_en = dataArray_57_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_7_cachedata_MPORT_addr = dataArray_57_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_7_cachedata_MPORT_data = dataArray_57_7[dataArray_57_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_7_MPORT_addr = replace_set;
  assign dataArray_57_7_MPORT_mask = _GEN_9008 & _GEN_7199;
  assign dataArray_57_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_8_cachedata_MPORT_en = dataArray_57_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_8_cachedata_MPORT_addr = dataArray_57_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_8_cachedata_MPORT_data = dataArray_57_8[dataArray_57_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_8_MPORT_addr = replace_set;
  assign dataArray_57_8_MPORT_mask = _GEN_9008 & _GEN_7201;
  assign dataArray_57_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_9_cachedata_MPORT_en = dataArray_57_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_9_cachedata_MPORT_addr = dataArray_57_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_9_cachedata_MPORT_data = dataArray_57_9[dataArray_57_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_9_MPORT_addr = replace_set;
  assign dataArray_57_9_MPORT_mask = _GEN_9008 & _GEN_7203;
  assign dataArray_57_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_10_cachedata_MPORT_en = dataArray_57_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_10_cachedata_MPORT_addr = dataArray_57_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_10_cachedata_MPORT_data = dataArray_57_10[dataArray_57_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_10_MPORT_addr = replace_set;
  assign dataArray_57_10_MPORT_mask = _GEN_9008 & _GEN_7205;
  assign dataArray_57_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_11_cachedata_MPORT_en = dataArray_57_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_11_cachedata_MPORT_addr = dataArray_57_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_11_cachedata_MPORT_data = dataArray_57_11[dataArray_57_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_11_MPORT_addr = replace_set;
  assign dataArray_57_11_MPORT_mask = _GEN_9008 & _GEN_7207;
  assign dataArray_57_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_12_cachedata_MPORT_en = dataArray_57_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_12_cachedata_MPORT_addr = dataArray_57_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_12_cachedata_MPORT_data = dataArray_57_12[dataArray_57_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_12_MPORT_addr = replace_set;
  assign dataArray_57_12_MPORT_mask = _GEN_9008 & _GEN_7209;
  assign dataArray_57_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_13_cachedata_MPORT_en = dataArray_57_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_13_cachedata_MPORT_addr = dataArray_57_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_13_cachedata_MPORT_data = dataArray_57_13[dataArray_57_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_13_MPORT_addr = replace_set;
  assign dataArray_57_13_MPORT_mask = _GEN_9008 & _GEN_7211;
  assign dataArray_57_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_14_cachedata_MPORT_en = dataArray_57_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_14_cachedata_MPORT_addr = dataArray_57_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_14_cachedata_MPORT_data = dataArray_57_14[dataArray_57_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_14_MPORT_addr = replace_set;
  assign dataArray_57_14_MPORT_mask = _GEN_9008 & _GEN_7213;
  assign dataArray_57_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_57_15_cachedata_MPORT_en = dataArray_57_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_57_15_cachedata_MPORT_addr = dataArray_57_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_57_15_cachedata_MPORT_data = dataArray_57_15[dataArray_57_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_57_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_57_15_MPORT_addr = replace_set;
  assign dataArray_57_15_MPORT_mask = _GEN_9008 & _GEN_7215;
  assign dataArray_57_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_0_cachedata_MPORT_en = dataArray_58_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_0_cachedata_MPORT_addr = dataArray_58_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_0_cachedata_MPORT_data = dataArray_58_0[dataArray_58_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_0_MPORT_addr = replace_set;
  assign dataArray_58_0_MPORT_mask = _GEN_9040 & _GEN_7185;
  assign dataArray_58_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_1_cachedata_MPORT_en = dataArray_58_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_1_cachedata_MPORT_addr = dataArray_58_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_1_cachedata_MPORT_data = dataArray_58_1[dataArray_58_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_1_MPORT_addr = replace_set;
  assign dataArray_58_1_MPORT_mask = _GEN_9040 & _GEN_7187;
  assign dataArray_58_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_2_cachedata_MPORT_en = dataArray_58_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_2_cachedata_MPORT_addr = dataArray_58_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_2_cachedata_MPORT_data = dataArray_58_2[dataArray_58_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_2_MPORT_addr = replace_set;
  assign dataArray_58_2_MPORT_mask = _GEN_9040 & _GEN_7189;
  assign dataArray_58_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_3_cachedata_MPORT_en = dataArray_58_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_3_cachedata_MPORT_addr = dataArray_58_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_3_cachedata_MPORT_data = dataArray_58_3[dataArray_58_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_3_MPORT_addr = replace_set;
  assign dataArray_58_3_MPORT_mask = _GEN_9040 & _GEN_7191;
  assign dataArray_58_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_4_cachedata_MPORT_en = dataArray_58_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_4_cachedata_MPORT_addr = dataArray_58_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_4_cachedata_MPORT_data = dataArray_58_4[dataArray_58_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_4_MPORT_addr = replace_set;
  assign dataArray_58_4_MPORT_mask = _GEN_9040 & _GEN_7193;
  assign dataArray_58_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_5_cachedata_MPORT_en = dataArray_58_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_5_cachedata_MPORT_addr = dataArray_58_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_5_cachedata_MPORT_data = dataArray_58_5[dataArray_58_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_5_MPORT_addr = replace_set;
  assign dataArray_58_5_MPORT_mask = _GEN_9040 & _GEN_7195;
  assign dataArray_58_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_6_cachedata_MPORT_en = dataArray_58_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_6_cachedata_MPORT_addr = dataArray_58_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_6_cachedata_MPORT_data = dataArray_58_6[dataArray_58_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_6_MPORT_addr = replace_set;
  assign dataArray_58_6_MPORT_mask = _GEN_9040 & _GEN_7197;
  assign dataArray_58_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_7_cachedata_MPORT_en = dataArray_58_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_7_cachedata_MPORT_addr = dataArray_58_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_7_cachedata_MPORT_data = dataArray_58_7[dataArray_58_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_7_MPORT_addr = replace_set;
  assign dataArray_58_7_MPORT_mask = _GEN_9040 & _GEN_7199;
  assign dataArray_58_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_8_cachedata_MPORT_en = dataArray_58_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_8_cachedata_MPORT_addr = dataArray_58_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_8_cachedata_MPORT_data = dataArray_58_8[dataArray_58_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_8_MPORT_addr = replace_set;
  assign dataArray_58_8_MPORT_mask = _GEN_9040 & _GEN_7201;
  assign dataArray_58_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_9_cachedata_MPORT_en = dataArray_58_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_9_cachedata_MPORT_addr = dataArray_58_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_9_cachedata_MPORT_data = dataArray_58_9[dataArray_58_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_9_MPORT_addr = replace_set;
  assign dataArray_58_9_MPORT_mask = _GEN_9040 & _GEN_7203;
  assign dataArray_58_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_10_cachedata_MPORT_en = dataArray_58_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_10_cachedata_MPORT_addr = dataArray_58_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_10_cachedata_MPORT_data = dataArray_58_10[dataArray_58_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_10_MPORT_addr = replace_set;
  assign dataArray_58_10_MPORT_mask = _GEN_9040 & _GEN_7205;
  assign dataArray_58_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_11_cachedata_MPORT_en = dataArray_58_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_11_cachedata_MPORT_addr = dataArray_58_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_11_cachedata_MPORT_data = dataArray_58_11[dataArray_58_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_11_MPORT_addr = replace_set;
  assign dataArray_58_11_MPORT_mask = _GEN_9040 & _GEN_7207;
  assign dataArray_58_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_12_cachedata_MPORT_en = dataArray_58_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_12_cachedata_MPORT_addr = dataArray_58_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_12_cachedata_MPORT_data = dataArray_58_12[dataArray_58_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_12_MPORT_addr = replace_set;
  assign dataArray_58_12_MPORT_mask = _GEN_9040 & _GEN_7209;
  assign dataArray_58_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_13_cachedata_MPORT_en = dataArray_58_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_13_cachedata_MPORT_addr = dataArray_58_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_13_cachedata_MPORT_data = dataArray_58_13[dataArray_58_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_13_MPORT_addr = replace_set;
  assign dataArray_58_13_MPORT_mask = _GEN_9040 & _GEN_7211;
  assign dataArray_58_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_14_cachedata_MPORT_en = dataArray_58_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_14_cachedata_MPORT_addr = dataArray_58_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_14_cachedata_MPORT_data = dataArray_58_14[dataArray_58_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_14_MPORT_addr = replace_set;
  assign dataArray_58_14_MPORT_mask = _GEN_9040 & _GEN_7213;
  assign dataArray_58_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_58_15_cachedata_MPORT_en = dataArray_58_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_58_15_cachedata_MPORT_addr = dataArray_58_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_58_15_cachedata_MPORT_data = dataArray_58_15[dataArray_58_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_58_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_58_15_MPORT_addr = replace_set;
  assign dataArray_58_15_MPORT_mask = _GEN_9040 & _GEN_7215;
  assign dataArray_58_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_0_cachedata_MPORT_en = dataArray_59_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_0_cachedata_MPORT_addr = dataArray_59_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_0_cachedata_MPORT_data = dataArray_59_0[dataArray_59_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_0_MPORT_addr = replace_set;
  assign dataArray_59_0_MPORT_mask = _GEN_9072 & _GEN_7185;
  assign dataArray_59_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_1_cachedata_MPORT_en = dataArray_59_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_1_cachedata_MPORT_addr = dataArray_59_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_1_cachedata_MPORT_data = dataArray_59_1[dataArray_59_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_1_MPORT_addr = replace_set;
  assign dataArray_59_1_MPORT_mask = _GEN_9072 & _GEN_7187;
  assign dataArray_59_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_2_cachedata_MPORT_en = dataArray_59_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_2_cachedata_MPORT_addr = dataArray_59_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_2_cachedata_MPORT_data = dataArray_59_2[dataArray_59_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_2_MPORT_addr = replace_set;
  assign dataArray_59_2_MPORT_mask = _GEN_9072 & _GEN_7189;
  assign dataArray_59_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_3_cachedata_MPORT_en = dataArray_59_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_3_cachedata_MPORT_addr = dataArray_59_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_3_cachedata_MPORT_data = dataArray_59_3[dataArray_59_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_3_MPORT_addr = replace_set;
  assign dataArray_59_3_MPORT_mask = _GEN_9072 & _GEN_7191;
  assign dataArray_59_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_4_cachedata_MPORT_en = dataArray_59_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_4_cachedata_MPORT_addr = dataArray_59_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_4_cachedata_MPORT_data = dataArray_59_4[dataArray_59_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_4_MPORT_addr = replace_set;
  assign dataArray_59_4_MPORT_mask = _GEN_9072 & _GEN_7193;
  assign dataArray_59_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_5_cachedata_MPORT_en = dataArray_59_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_5_cachedata_MPORT_addr = dataArray_59_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_5_cachedata_MPORT_data = dataArray_59_5[dataArray_59_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_5_MPORT_addr = replace_set;
  assign dataArray_59_5_MPORT_mask = _GEN_9072 & _GEN_7195;
  assign dataArray_59_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_6_cachedata_MPORT_en = dataArray_59_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_6_cachedata_MPORT_addr = dataArray_59_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_6_cachedata_MPORT_data = dataArray_59_6[dataArray_59_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_6_MPORT_addr = replace_set;
  assign dataArray_59_6_MPORT_mask = _GEN_9072 & _GEN_7197;
  assign dataArray_59_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_7_cachedata_MPORT_en = dataArray_59_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_7_cachedata_MPORT_addr = dataArray_59_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_7_cachedata_MPORT_data = dataArray_59_7[dataArray_59_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_7_MPORT_addr = replace_set;
  assign dataArray_59_7_MPORT_mask = _GEN_9072 & _GEN_7199;
  assign dataArray_59_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_8_cachedata_MPORT_en = dataArray_59_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_8_cachedata_MPORT_addr = dataArray_59_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_8_cachedata_MPORT_data = dataArray_59_8[dataArray_59_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_8_MPORT_addr = replace_set;
  assign dataArray_59_8_MPORT_mask = _GEN_9072 & _GEN_7201;
  assign dataArray_59_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_9_cachedata_MPORT_en = dataArray_59_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_9_cachedata_MPORT_addr = dataArray_59_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_9_cachedata_MPORT_data = dataArray_59_9[dataArray_59_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_9_MPORT_addr = replace_set;
  assign dataArray_59_9_MPORT_mask = _GEN_9072 & _GEN_7203;
  assign dataArray_59_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_10_cachedata_MPORT_en = dataArray_59_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_10_cachedata_MPORT_addr = dataArray_59_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_10_cachedata_MPORT_data = dataArray_59_10[dataArray_59_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_10_MPORT_addr = replace_set;
  assign dataArray_59_10_MPORT_mask = _GEN_9072 & _GEN_7205;
  assign dataArray_59_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_11_cachedata_MPORT_en = dataArray_59_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_11_cachedata_MPORT_addr = dataArray_59_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_11_cachedata_MPORT_data = dataArray_59_11[dataArray_59_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_11_MPORT_addr = replace_set;
  assign dataArray_59_11_MPORT_mask = _GEN_9072 & _GEN_7207;
  assign dataArray_59_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_12_cachedata_MPORT_en = dataArray_59_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_12_cachedata_MPORT_addr = dataArray_59_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_12_cachedata_MPORT_data = dataArray_59_12[dataArray_59_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_12_MPORT_addr = replace_set;
  assign dataArray_59_12_MPORT_mask = _GEN_9072 & _GEN_7209;
  assign dataArray_59_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_13_cachedata_MPORT_en = dataArray_59_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_13_cachedata_MPORT_addr = dataArray_59_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_13_cachedata_MPORT_data = dataArray_59_13[dataArray_59_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_13_MPORT_addr = replace_set;
  assign dataArray_59_13_MPORT_mask = _GEN_9072 & _GEN_7211;
  assign dataArray_59_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_14_cachedata_MPORT_en = dataArray_59_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_14_cachedata_MPORT_addr = dataArray_59_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_14_cachedata_MPORT_data = dataArray_59_14[dataArray_59_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_14_MPORT_addr = replace_set;
  assign dataArray_59_14_MPORT_mask = _GEN_9072 & _GEN_7213;
  assign dataArray_59_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_59_15_cachedata_MPORT_en = dataArray_59_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_59_15_cachedata_MPORT_addr = dataArray_59_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_59_15_cachedata_MPORT_data = dataArray_59_15[dataArray_59_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_59_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_59_15_MPORT_addr = replace_set;
  assign dataArray_59_15_MPORT_mask = _GEN_9072 & _GEN_7215;
  assign dataArray_59_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_0_cachedata_MPORT_en = dataArray_60_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_0_cachedata_MPORT_addr = dataArray_60_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_0_cachedata_MPORT_data = dataArray_60_0[dataArray_60_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_0_MPORT_addr = replace_set;
  assign dataArray_60_0_MPORT_mask = _GEN_9104 & _GEN_7185;
  assign dataArray_60_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_1_cachedata_MPORT_en = dataArray_60_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_1_cachedata_MPORT_addr = dataArray_60_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_1_cachedata_MPORT_data = dataArray_60_1[dataArray_60_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_1_MPORT_addr = replace_set;
  assign dataArray_60_1_MPORT_mask = _GEN_9104 & _GEN_7187;
  assign dataArray_60_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_2_cachedata_MPORT_en = dataArray_60_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_2_cachedata_MPORT_addr = dataArray_60_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_2_cachedata_MPORT_data = dataArray_60_2[dataArray_60_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_2_MPORT_addr = replace_set;
  assign dataArray_60_2_MPORT_mask = _GEN_9104 & _GEN_7189;
  assign dataArray_60_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_3_cachedata_MPORT_en = dataArray_60_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_3_cachedata_MPORT_addr = dataArray_60_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_3_cachedata_MPORT_data = dataArray_60_3[dataArray_60_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_3_MPORT_addr = replace_set;
  assign dataArray_60_3_MPORT_mask = _GEN_9104 & _GEN_7191;
  assign dataArray_60_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_4_cachedata_MPORT_en = dataArray_60_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_4_cachedata_MPORT_addr = dataArray_60_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_4_cachedata_MPORT_data = dataArray_60_4[dataArray_60_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_4_MPORT_addr = replace_set;
  assign dataArray_60_4_MPORT_mask = _GEN_9104 & _GEN_7193;
  assign dataArray_60_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_5_cachedata_MPORT_en = dataArray_60_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_5_cachedata_MPORT_addr = dataArray_60_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_5_cachedata_MPORT_data = dataArray_60_5[dataArray_60_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_5_MPORT_addr = replace_set;
  assign dataArray_60_5_MPORT_mask = _GEN_9104 & _GEN_7195;
  assign dataArray_60_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_6_cachedata_MPORT_en = dataArray_60_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_6_cachedata_MPORT_addr = dataArray_60_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_6_cachedata_MPORT_data = dataArray_60_6[dataArray_60_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_6_MPORT_addr = replace_set;
  assign dataArray_60_6_MPORT_mask = _GEN_9104 & _GEN_7197;
  assign dataArray_60_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_7_cachedata_MPORT_en = dataArray_60_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_7_cachedata_MPORT_addr = dataArray_60_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_7_cachedata_MPORT_data = dataArray_60_7[dataArray_60_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_7_MPORT_addr = replace_set;
  assign dataArray_60_7_MPORT_mask = _GEN_9104 & _GEN_7199;
  assign dataArray_60_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_8_cachedata_MPORT_en = dataArray_60_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_8_cachedata_MPORT_addr = dataArray_60_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_8_cachedata_MPORT_data = dataArray_60_8[dataArray_60_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_8_MPORT_addr = replace_set;
  assign dataArray_60_8_MPORT_mask = _GEN_9104 & _GEN_7201;
  assign dataArray_60_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_9_cachedata_MPORT_en = dataArray_60_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_9_cachedata_MPORT_addr = dataArray_60_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_9_cachedata_MPORT_data = dataArray_60_9[dataArray_60_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_9_MPORT_addr = replace_set;
  assign dataArray_60_9_MPORT_mask = _GEN_9104 & _GEN_7203;
  assign dataArray_60_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_10_cachedata_MPORT_en = dataArray_60_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_10_cachedata_MPORT_addr = dataArray_60_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_10_cachedata_MPORT_data = dataArray_60_10[dataArray_60_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_10_MPORT_addr = replace_set;
  assign dataArray_60_10_MPORT_mask = _GEN_9104 & _GEN_7205;
  assign dataArray_60_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_11_cachedata_MPORT_en = dataArray_60_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_11_cachedata_MPORT_addr = dataArray_60_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_11_cachedata_MPORT_data = dataArray_60_11[dataArray_60_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_11_MPORT_addr = replace_set;
  assign dataArray_60_11_MPORT_mask = _GEN_9104 & _GEN_7207;
  assign dataArray_60_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_12_cachedata_MPORT_en = dataArray_60_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_12_cachedata_MPORT_addr = dataArray_60_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_12_cachedata_MPORT_data = dataArray_60_12[dataArray_60_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_12_MPORT_addr = replace_set;
  assign dataArray_60_12_MPORT_mask = _GEN_9104 & _GEN_7209;
  assign dataArray_60_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_13_cachedata_MPORT_en = dataArray_60_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_13_cachedata_MPORT_addr = dataArray_60_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_13_cachedata_MPORT_data = dataArray_60_13[dataArray_60_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_13_MPORT_addr = replace_set;
  assign dataArray_60_13_MPORT_mask = _GEN_9104 & _GEN_7211;
  assign dataArray_60_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_14_cachedata_MPORT_en = dataArray_60_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_14_cachedata_MPORT_addr = dataArray_60_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_14_cachedata_MPORT_data = dataArray_60_14[dataArray_60_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_14_MPORT_addr = replace_set;
  assign dataArray_60_14_MPORT_mask = _GEN_9104 & _GEN_7213;
  assign dataArray_60_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_60_15_cachedata_MPORT_en = dataArray_60_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_60_15_cachedata_MPORT_addr = dataArray_60_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_60_15_cachedata_MPORT_data = dataArray_60_15[dataArray_60_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_60_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_60_15_MPORT_addr = replace_set;
  assign dataArray_60_15_MPORT_mask = _GEN_9104 & _GEN_7215;
  assign dataArray_60_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_0_cachedata_MPORT_en = dataArray_61_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_0_cachedata_MPORT_addr = dataArray_61_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_0_cachedata_MPORT_data = dataArray_61_0[dataArray_61_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_0_MPORT_addr = replace_set;
  assign dataArray_61_0_MPORT_mask = _GEN_9136 & _GEN_7185;
  assign dataArray_61_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_1_cachedata_MPORT_en = dataArray_61_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_1_cachedata_MPORT_addr = dataArray_61_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_1_cachedata_MPORT_data = dataArray_61_1[dataArray_61_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_1_MPORT_addr = replace_set;
  assign dataArray_61_1_MPORT_mask = _GEN_9136 & _GEN_7187;
  assign dataArray_61_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_2_cachedata_MPORT_en = dataArray_61_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_2_cachedata_MPORT_addr = dataArray_61_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_2_cachedata_MPORT_data = dataArray_61_2[dataArray_61_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_2_MPORT_addr = replace_set;
  assign dataArray_61_2_MPORT_mask = _GEN_9136 & _GEN_7189;
  assign dataArray_61_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_3_cachedata_MPORT_en = dataArray_61_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_3_cachedata_MPORT_addr = dataArray_61_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_3_cachedata_MPORT_data = dataArray_61_3[dataArray_61_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_3_MPORT_addr = replace_set;
  assign dataArray_61_3_MPORT_mask = _GEN_9136 & _GEN_7191;
  assign dataArray_61_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_4_cachedata_MPORT_en = dataArray_61_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_4_cachedata_MPORT_addr = dataArray_61_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_4_cachedata_MPORT_data = dataArray_61_4[dataArray_61_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_4_MPORT_addr = replace_set;
  assign dataArray_61_4_MPORT_mask = _GEN_9136 & _GEN_7193;
  assign dataArray_61_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_5_cachedata_MPORT_en = dataArray_61_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_5_cachedata_MPORT_addr = dataArray_61_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_5_cachedata_MPORT_data = dataArray_61_5[dataArray_61_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_5_MPORT_addr = replace_set;
  assign dataArray_61_5_MPORT_mask = _GEN_9136 & _GEN_7195;
  assign dataArray_61_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_6_cachedata_MPORT_en = dataArray_61_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_6_cachedata_MPORT_addr = dataArray_61_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_6_cachedata_MPORT_data = dataArray_61_6[dataArray_61_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_6_MPORT_addr = replace_set;
  assign dataArray_61_6_MPORT_mask = _GEN_9136 & _GEN_7197;
  assign dataArray_61_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_7_cachedata_MPORT_en = dataArray_61_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_7_cachedata_MPORT_addr = dataArray_61_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_7_cachedata_MPORT_data = dataArray_61_7[dataArray_61_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_7_MPORT_addr = replace_set;
  assign dataArray_61_7_MPORT_mask = _GEN_9136 & _GEN_7199;
  assign dataArray_61_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_8_cachedata_MPORT_en = dataArray_61_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_8_cachedata_MPORT_addr = dataArray_61_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_8_cachedata_MPORT_data = dataArray_61_8[dataArray_61_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_8_MPORT_addr = replace_set;
  assign dataArray_61_8_MPORT_mask = _GEN_9136 & _GEN_7201;
  assign dataArray_61_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_9_cachedata_MPORT_en = dataArray_61_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_9_cachedata_MPORT_addr = dataArray_61_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_9_cachedata_MPORT_data = dataArray_61_9[dataArray_61_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_9_MPORT_addr = replace_set;
  assign dataArray_61_9_MPORT_mask = _GEN_9136 & _GEN_7203;
  assign dataArray_61_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_10_cachedata_MPORT_en = dataArray_61_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_10_cachedata_MPORT_addr = dataArray_61_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_10_cachedata_MPORT_data = dataArray_61_10[dataArray_61_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_10_MPORT_addr = replace_set;
  assign dataArray_61_10_MPORT_mask = _GEN_9136 & _GEN_7205;
  assign dataArray_61_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_11_cachedata_MPORT_en = dataArray_61_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_11_cachedata_MPORT_addr = dataArray_61_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_11_cachedata_MPORT_data = dataArray_61_11[dataArray_61_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_11_MPORT_addr = replace_set;
  assign dataArray_61_11_MPORT_mask = _GEN_9136 & _GEN_7207;
  assign dataArray_61_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_12_cachedata_MPORT_en = dataArray_61_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_12_cachedata_MPORT_addr = dataArray_61_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_12_cachedata_MPORT_data = dataArray_61_12[dataArray_61_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_12_MPORT_addr = replace_set;
  assign dataArray_61_12_MPORT_mask = _GEN_9136 & _GEN_7209;
  assign dataArray_61_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_13_cachedata_MPORT_en = dataArray_61_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_13_cachedata_MPORT_addr = dataArray_61_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_13_cachedata_MPORT_data = dataArray_61_13[dataArray_61_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_13_MPORT_addr = replace_set;
  assign dataArray_61_13_MPORT_mask = _GEN_9136 & _GEN_7211;
  assign dataArray_61_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_14_cachedata_MPORT_en = dataArray_61_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_14_cachedata_MPORT_addr = dataArray_61_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_14_cachedata_MPORT_data = dataArray_61_14[dataArray_61_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_14_MPORT_addr = replace_set;
  assign dataArray_61_14_MPORT_mask = _GEN_9136 & _GEN_7213;
  assign dataArray_61_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_61_15_cachedata_MPORT_en = dataArray_61_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_61_15_cachedata_MPORT_addr = dataArray_61_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_61_15_cachedata_MPORT_data = dataArray_61_15[dataArray_61_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_61_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_61_15_MPORT_addr = replace_set;
  assign dataArray_61_15_MPORT_mask = _GEN_9136 & _GEN_7215;
  assign dataArray_61_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_0_cachedata_MPORT_en = dataArray_62_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_0_cachedata_MPORT_addr = dataArray_62_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_0_cachedata_MPORT_data = dataArray_62_0[dataArray_62_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_0_MPORT_addr = replace_set;
  assign dataArray_62_0_MPORT_mask = _GEN_9168 & _GEN_7185;
  assign dataArray_62_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_1_cachedata_MPORT_en = dataArray_62_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_1_cachedata_MPORT_addr = dataArray_62_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_1_cachedata_MPORT_data = dataArray_62_1[dataArray_62_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_1_MPORT_addr = replace_set;
  assign dataArray_62_1_MPORT_mask = _GEN_9168 & _GEN_7187;
  assign dataArray_62_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_2_cachedata_MPORT_en = dataArray_62_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_2_cachedata_MPORT_addr = dataArray_62_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_2_cachedata_MPORT_data = dataArray_62_2[dataArray_62_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_2_MPORT_addr = replace_set;
  assign dataArray_62_2_MPORT_mask = _GEN_9168 & _GEN_7189;
  assign dataArray_62_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_3_cachedata_MPORT_en = dataArray_62_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_3_cachedata_MPORT_addr = dataArray_62_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_3_cachedata_MPORT_data = dataArray_62_3[dataArray_62_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_3_MPORT_addr = replace_set;
  assign dataArray_62_3_MPORT_mask = _GEN_9168 & _GEN_7191;
  assign dataArray_62_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_4_cachedata_MPORT_en = dataArray_62_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_4_cachedata_MPORT_addr = dataArray_62_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_4_cachedata_MPORT_data = dataArray_62_4[dataArray_62_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_4_MPORT_addr = replace_set;
  assign dataArray_62_4_MPORT_mask = _GEN_9168 & _GEN_7193;
  assign dataArray_62_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_5_cachedata_MPORT_en = dataArray_62_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_5_cachedata_MPORT_addr = dataArray_62_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_5_cachedata_MPORT_data = dataArray_62_5[dataArray_62_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_5_MPORT_addr = replace_set;
  assign dataArray_62_5_MPORT_mask = _GEN_9168 & _GEN_7195;
  assign dataArray_62_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_6_cachedata_MPORT_en = dataArray_62_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_6_cachedata_MPORT_addr = dataArray_62_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_6_cachedata_MPORT_data = dataArray_62_6[dataArray_62_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_6_MPORT_addr = replace_set;
  assign dataArray_62_6_MPORT_mask = _GEN_9168 & _GEN_7197;
  assign dataArray_62_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_7_cachedata_MPORT_en = dataArray_62_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_7_cachedata_MPORT_addr = dataArray_62_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_7_cachedata_MPORT_data = dataArray_62_7[dataArray_62_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_7_MPORT_addr = replace_set;
  assign dataArray_62_7_MPORT_mask = _GEN_9168 & _GEN_7199;
  assign dataArray_62_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_8_cachedata_MPORT_en = dataArray_62_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_8_cachedata_MPORT_addr = dataArray_62_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_8_cachedata_MPORT_data = dataArray_62_8[dataArray_62_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_8_MPORT_addr = replace_set;
  assign dataArray_62_8_MPORT_mask = _GEN_9168 & _GEN_7201;
  assign dataArray_62_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_9_cachedata_MPORT_en = dataArray_62_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_9_cachedata_MPORT_addr = dataArray_62_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_9_cachedata_MPORT_data = dataArray_62_9[dataArray_62_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_9_MPORT_addr = replace_set;
  assign dataArray_62_9_MPORT_mask = _GEN_9168 & _GEN_7203;
  assign dataArray_62_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_10_cachedata_MPORT_en = dataArray_62_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_10_cachedata_MPORT_addr = dataArray_62_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_10_cachedata_MPORT_data = dataArray_62_10[dataArray_62_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_10_MPORT_addr = replace_set;
  assign dataArray_62_10_MPORT_mask = _GEN_9168 & _GEN_7205;
  assign dataArray_62_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_11_cachedata_MPORT_en = dataArray_62_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_11_cachedata_MPORT_addr = dataArray_62_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_11_cachedata_MPORT_data = dataArray_62_11[dataArray_62_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_11_MPORT_addr = replace_set;
  assign dataArray_62_11_MPORT_mask = _GEN_9168 & _GEN_7207;
  assign dataArray_62_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_12_cachedata_MPORT_en = dataArray_62_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_12_cachedata_MPORT_addr = dataArray_62_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_12_cachedata_MPORT_data = dataArray_62_12[dataArray_62_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_12_MPORT_addr = replace_set;
  assign dataArray_62_12_MPORT_mask = _GEN_9168 & _GEN_7209;
  assign dataArray_62_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_13_cachedata_MPORT_en = dataArray_62_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_13_cachedata_MPORT_addr = dataArray_62_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_13_cachedata_MPORT_data = dataArray_62_13[dataArray_62_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_13_MPORT_addr = replace_set;
  assign dataArray_62_13_MPORT_mask = _GEN_9168 & _GEN_7211;
  assign dataArray_62_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_14_cachedata_MPORT_en = dataArray_62_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_14_cachedata_MPORT_addr = dataArray_62_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_14_cachedata_MPORT_data = dataArray_62_14[dataArray_62_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_14_MPORT_addr = replace_set;
  assign dataArray_62_14_MPORT_mask = _GEN_9168 & _GEN_7213;
  assign dataArray_62_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_62_15_cachedata_MPORT_en = dataArray_62_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_62_15_cachedata_MPORT_addr = dataArray_62_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_62_15_cachedata_MPORT_data = dataArray_62_15[dataArray_62_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_62_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_62_15_MPORT_addr = replace_set;
  assign dataArray_62_15_MPORT_mask = _GEN_9168 & _GEN_7215;
  assign dataArray_62_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_0_cachedata_MPORT_en = dataArray_63_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_0_cachedata_MPORT_addr = dataArray_63_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_0_cachedata_MPORT_data = dataArray_63_0[dataArray_63_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_0_MPORT_addr = replace_set;
  assign dataArray_63_0_MPORT_mask = _GEN_9200 & _GEN_7185;
  assign dataArray_63_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_1_cachedata_MPORT_en = dataArray_63_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_1_cachedata_MPORT_addr = dataArray_63_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_1_cachedata_MPORT_data = dataArray_63_1[dataArray_63_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_1_MPORT_addr = replace_set;
  assign dataArray_63_1_MPORT_mask = _GEN_9200 & _GEN_7187;
  assign dataArray_63_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_2_cachedata_MPORT_en = dataArray_63_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_2_cachedata_MPORT_addr = dataArray_63_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_2_cachedata_MPORT_data = dataArray_63_2[dataArray_63_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_2_MPORT_addr = replace_set;
  assign dataArray_63_2_MPORT_mask = _GEN_9200 & _GEN_7189;
  assign dataArray_63_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_3_cachedata_MPORT_en = dataArray_63_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_3_cachedata_MPORT_addr = dataArray_63_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_3_cachedata_MPORT_data = dataArray_63_3[dataArray_63_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_3_MPORT_addr = replace_set;
  assign dataArray_63_3_MPORT_mask = _GEN_9200 & _GEN_7191;
  assign dataArray_63_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_4_cachedata_MPORT_en = dataArray_63_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_4_cachedata_MPORT_addr = dataArray_63_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_4_cachedata_MPORT_data = dataArray_63_4[dataArray_63_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_4_MPORT_addr = replace_set;
  assign dataArray_63_4_MPORT_mask = _GEN_9200 & _GEN_7193;
  assign dataArray_63_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_5_cachedata_MPORT_en = dataArray_63_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_5_cachedata_MPORT_addr = dataArray_63_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_5_cachedata_MPORT_data = dataArray_63_5[dataArray_63_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_5_MPORT_addr = replace_set;
  assign dataArray_63_5_MPORT_mask = _GEN_9200 & _GEN_7195;
  assign dataArray_63_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_6_cachedata_MPORT_en = dataArray_63_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_6_cachedata_MPORT_addr = dataArray_63_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_6_cachedata_MPORT_data = dataArray_63_6[dataArray_63_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_6_MPORT_addr = replace_set;
  assign dataArray_63_6_MPORT_mask = _GEN_9200 & _GEN_7197;
  assign dataArray_63_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_7_cachedata_MPORT_en = dataArray_63_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_7_cachedata_MPORT_addr = dataArray_63_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_7_cachedata_MPORT_data = dataArray_63_7[dataArray_63_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_7_MPORT_addr = replace_set;
  assign dataArray_63_7_MPORT_mask = _GEN_9200 & _GEN_7199;
  assign dataArray_63_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_8_cachedata_MPORT_en = dataArray_63_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_8_cachedata_MPORT_addr = dataArray_63_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_8_cachedata_MPORT_data = dataArray_63_8[dataArray_63_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_8_MPORT_addr = replace_set;
  assign dataArray_63_8_MPORT_mask = _GEN_9200 & _GEN_7201;
  assign dataArray_63_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_9_cachedata_MPORT_en = dataArray_63_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_9_cachedata_MPORT_addr = dataArray_63_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_9_cachedata_MPORT_data = dataArray_63_9[dataArray_63_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_9_MPORT_addr = replace_set;
  assign dataArray_63_9_MPORT_mask = _GEN_9200 & _GEN_7203;
  assign dataArray_63_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_10_cachedata_MPORT_en = dataArray_63_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_10_cachedata_MPORT_addr = dataArray_63_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_10_cachedata_MPORT_data = dataArray_63_10[dataArray_63_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_10_MPORT_addr = replace_set;
  assign dataArray_63_10_MPORT_mask = _GEN_9200 & _GEN_7205;
  assign dataArray_63_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_11_cachedata_MPORT_en = dataArray_63_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_11_cachedata_MPORT_addr = dataArray_63_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_11_cachedata_MPORT_data = dataArray_63_11[dataArray_63_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_11_MPORT_addr = replace_set;
  assign dataArray_63_11_MPORT_mask = _GEN_9200 & _GEN_7207;
  assign dataArray_63_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_12_cachedata_MPORT_en = dataArray_63_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_12_cachedata_MPORT_addr = dataArray_63_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_12_cachedata_MPORT_data = dataArray_63_12[dataArray_63_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_12_MPORT_addr = replace_set;
  assign dataArray_63_12_MPORT_mask = _GEN_9200 & _GEN_7209;
  assign dataArray_63_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_13_cachedata_MPORT_en = dataArray_63_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_13_cachedata_MPORT_addr = dataArray_63_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_13_cachedata_MPORT_data = dataArray_63_13[dataArray_63_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_13_MPORT_addr = replace_set;
  assign dataArray_63_13_MPORT_mask = _GEN_9200 & _GEN_7211;
  assign dataArray_63_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_14_cachedata_MPORT_en = dataArray_63_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_14_cachedata_MPORT_addr = dataArray_63_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_14_cachedata_MPORT_data = dataArray_63_14[dataArray_63_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_14_MPORT_addr = replace_set;
  assign dataArray_63_14_MPORT_mask = _GEN_9200 & _GEN_7213;
  assign dataArray_63_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_63_15_cachedata_MPORT_en = dataArray_63_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_63_15_cachedata_MPORT_addr = dataArray_63_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_63_15_cachedata_MPORT_data = dataArray_63_15[dataArray_63_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_63_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_63_15_MPORT_addr = replace_set;
  assign dataArray_63_15_MPORT_mask = _GEN_9200 & _GEN_7215;
  assign dataArray_63_15_MPORT_en = _T_6 & _off_T;
  assign from_IFU_ready = 3'h0 == state_cache; // @[Mux.scala 81:61]
  assign to_IFU_valid = 3'h1 == state_cache; // @[Mux.scala 81:61]
  assign to_IFU_bits_data = hit ? _GEN_7183 : 32'h13; // @[cache.scala 108:28]
  assign to_sram_ar_valid = 3'h2 == state_cache; // @[Mux.scala 81:61]
  assign to_sram_ar_bits_addr = _to_sram_ar_bits_addr_T_3[31:0]; // @[cache.scala 91:27]
  assign to_sram_ar_bits_len = {{4'd0}, _to_sram_ar_bits_len_T_1}; // @[cache.scala 93:27]
  assign to_sram_r_ready = 3'h3 == state_cache; // @[Mux.scala 81:61]
  always @(posedge clock) begin
    if (dataArray_0_0_MPORT_en & dataArray_0_0_MPORT_mask) begin
      dataArray_0_0[dataArray_0_0_MPORT_addr] <= dataArray_0_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_1_MPORT_en & dataArray_0_1_MPORT_mask) begin
      dataArray_0_1[dataArray_0_1_MPORT_addr] <= dataArray_0_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_2_MPORT_en & dataArray_0_2_MPORT_mask) begin
      dataArray_0_2[dataArray_0_2_MPORT_addr] <= dataArray_0_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_3_MPORT_en & dataArray_0_3_MPORT_mask) begin
      dataArray_0_3[dataArray_0_3_MPORT_addr] <= dataArray_0_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_4_MPORT_en & dataArray_0_4_MPORT_mask) begin
      dataArray_0_4[dataArray_0_4_MPORT_addr] <= dataArray_0_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_5_MPORT_en & dataArray_0_5_MPORT_mask) begin
      dataArray_0_5[dataArray_0_5_MPORT_addr] <= dataArray_0_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_6_MPORT_en & dataArray_0_6_MPORT_mask) begin
      dataArray_0_6[dataArray_0_6_MPORT_addr] <= dataArray_0_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_7_MPORT_en & dataArray_0_7_MPORT_mask) begin
      dataArray_0_7[dataArray_0_7_MPORT_addr] <= dataArray_0_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_8_MPORT_en & dataArray_0_8_MPORT_mask) begin
      dataArray_0_8[dataArray_0_8_MPORT_addr] <= dataArray_0_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_9_MPORT_en & dataArray_0_9_MPORT_mask) begin
      dataArray_0_9[dataArray_0_9_MPORT_addr] <= dataArray_0_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_10_MPORT_en & dataArray_0_10_MPORT_mask) begin
      dataArray_0_10[dataArray_0_10_MPORT_addr] <= dataArray_0_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_11_MPORT_en & dataArray_0_11_MPORT_mask) begin
      dataArray_0_11[dataArray_0_11_MPORT_addr] <= dataArray_0_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_12_MPORT_en & dataArray_0_12_MPORT_mask) begin
      dataArray_0_12[dataArray_0_12_MPORT_addr] <= dataArray_0_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_13_MPORT_en & dataArray_0_13_MPORT_mask) begin
      dataArray_0_13[dataArray_0_13_MPORT_addr] <= dataArray_0_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_14_MPORT_en & dataArray_0_14_MPORT_mask) begin
      dataArray_0_14[dataArray_0_14_MPORT_addr] <= dataArray_0_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_0_15_MPORT_en & dataArray_0_15_MPORT_mask) begin
      dataArray_0_15[dataArray_0_15_MPORT_addr] <= dataArray_0_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_0_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_0_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_0_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_0_MPORT_en & dataArray_1_0_MPORT_mask) begin
      dataArray_1_0[dataArray_1_0_MPORT_addr] <= dataArray_1_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_1_MPORT_en & dataArray_1_1_MPORT_mask) begin
      dataArray_1_1[dataArray_1_1_MPORT_addr] <= dataArray_1_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_2_MPORT_en & dataArray_1_2_MPORT_mask) begin
      dataArray_1_2[dataArray_1_2_MPORT_addr] <= dataArray_1_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_3_MPORT_en & dataArray_1_3_MPORT_mask) begin
      dataArray_1_3[dataArray_1_3_MPORT_addr] <= dataArray_1_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_4_MPORT_en & dataArray_1_4_MPORT_mask) begin
      dataArray_1_4[dataArray_1_4_MPORT_addr] <= dataArray_1_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_5_MPORT_en & dataArray_1_5_MPORT_mask) begin
      dataArray_1_5[dataArray_1_5_MPORT_addr] <= dataArray_1_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_6_MPORT_en & dataArray_1_6_MPORT_mask) begin
      dataArray_1_6[dataArray_1_6_MPORT_addr] <= dataArray_1_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_7_MPORT_en & dataArray_1_7_MPORT_mask) begin
      dataArray_1_7[dataArray_1_7_MPORT_addr] <= dataArray_1_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_8_MPORT_en & dataArray_1_8_MPORT_mask) begin
      dataArray_1_8[dataArray_1_8_MPORT_addr] <= dataArray_1_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_9_MPORT_en & dataArray_1_9_MPORT_mask) begin
      dataArray_1_9[dataArray_1_9_MPORT_addr] <= dataArray_1_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_10_MPORT_en & dataArray_1_10_MPORT_mask) begin
      dataArray_1_10[dataArray_1_10_MPORT_addr] <= dataArray_1_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_11_MPORT_en & dataArray_1_11_MPORT_mask) begin
      dataArray_1_11[dataArray_1_11_MPORT_addr] <= dataArray_1_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_12_MPORT_en & dataArray_1_12_MPORT_mask) begin
      dataArray_1_12[dataArray_1_12_MPORT_addr] <= dataArray_1_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_13_MPORT_en & dataArray_1_13_MPORT_mask) begin
      dataArray_1_13[dataArray_1_13_MPORT_addr] <= dataArray_1_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_14_MPORT_en & dataArray_1_14_MPORT_mask) begin
      dataArray_1_14[dataArray_1_14_MPORT_addr] <= dataArray_1_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_1_15_MPORT_en & dataArray_1_15_MPORT_mask) begin
      dataArray_1_15[dataArray_1_15_MPORT_addr] <= dataArray_1_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_1_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_1_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_1_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_0_MPORT_en & dataArray_2_0_MPORT_mask) begin
      dataArray_2_0[dataArray_2_0_MPORT_addr] <= dataArray_2_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_1_MPORT_en & dataArray_2_1_MPORT_mask) begin
      dataArray_2_1[dataArray_2_1_MPORT_addr] <= dataArray_2_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_2_MPORT_en & dataArray_2_2_MPORT_mask) begin
      dataArray_2_2[dataArray_2_2_MPORT_addr] <= dataArray_2_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_3_MPORT_en & dataArray_2_3_MPORT_mask) begin
      dataArray_2_3[dataArray_2_3_MPORT_addr] <= dataArray_2_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_4_MPORT_en & dataArray_2_4_MPORT_mask) begin
      dataArray_2_4[dataArray_2_4_MPORT_addr] <= dataArray_2_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_5_MPORT_en & dataArray_2_5_MPORT_mask) begin
      dataArray_2_5[dataArray_2_5_MPORT_addr] <= dataArray_2_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_6_MPORT_en & dataArray_2_6_MPORT_mask) begin
      dataArray_2_6[dataArray_2_6_MPORT_addr] <= dataArray_2_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_7_MPORT_en & dataArray_2_7_MPORT_mask) begin
      dataArray_2_7[dataArray_2_7_MPORT_addr] <= dataArray_2_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_8_MPORT_en & dataArray_2_8_MPORT_mask) begin
      dataArray_2_8[dataArray_2_8_MPORT_addr] <= dataArray_2_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_9_MPORT_en & dataArray_2_9_MPORT_mask) begin
      dataArray_2_9[dataArray_2_9_MPORT_addr] <= dataArray_2_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_10_MPORT_en & dataArray_2_10_MPORT_mask) begin
      dataArray_2_10[dataArray_2_10_MPORT_addr] <= dataArray_2_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_11_MPORT_en & dataArray_2_11_MPORT_mask) begin
      dataArray_2_11[dataArray_2_11_MPORT_addr] <= dataArray_2_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_12_MPORT_en & dataArray_2_12_MPORT_mask) begin
      dataArray_2_12[dataArray_2_12_MPORT_addr] <= dataArray_2_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_13_MPORT_en & dataArray_2_13_MPORT_mask) begin
      dataArray_2_13[dataArray_2_13_MPORT_addr] <= dataArray_2_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_14_MPORT_en & dataArray_2_14_MPORT_mask) begin
      dataArray_2_14[dataArray_2_14_MPORT_addr] <= dataArray_2_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_2_15_MPORT_en & dataArray_2_15_MPORT_mask) begin
      dataArray_2_15[dataArray_2_15_MPORT_addr] <= dataArray_2_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_2_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_2_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_2_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_0_MPORT_en & dataArray_3_0_MPORT_mask) begin
      dataArray_3_0[dataArray_3_0_MPORT_addr] <= dataArray_3_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_1_MPORT_en & dataArray_3_1_MPORT_mask) begin
      dataArray_3_1[dataArray_3_1_MPORT_addr] <= dataArray_3_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_2_MPORT_en & dataArray_3_2_MPORT_mask) begin
      dataArray_3_2[dataArray_3_2_MPORT_addr] <= dataArray_3_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_3_MPORT_en & dataArray_3_3_MPORT_mask) begin
      dataArray_3_3[dataArray_3_3_MPORT_addr] <= dataArray_3_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_4_MPORT_en & dataArray_3_4_MPORT_mask) begin
      dataArray_3_4[dataArray_3_4_MPORT_addr] <= dataArray_3_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_5_MPORT_en & dataArray_3_5_MPORT_mask) begin
      dataArray_3_5[dataArray_3_5_MPORT_addr] <= dataArray_3_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_6_MPORT_en & dataArray_3_6_MPORT_mask) begin
      dataArray_3_6[dataArray_3_6_MPORT_addr] <= dataArray_3_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_7_MPORT_en & dataArray_3_7_MPORT_mask) begin
      dataArray_3_7[dataArray_3_7_MPORT_addr] <= dataArray_3_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_8_MPORT_en & dataArray_3_8_MPORT_mask) begin
      dataArray_3_8[dataArray_3_8_MPORT_addr] <= dataArray_3_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_9_MPORT_en & dataArray_3_9_MPORT_mask) begin
      dataArray_3_9[dataArray_3_9_MPORT_addr] <= dataArray_3_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_10_MPORT_en & dataArray_3_10_MPORT_mask) begin
      dataArray_3_10[dataArray_3_10_MPORT_addr] <= dataArray_3_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_11_MPORT_en & dataArray_3_11_MPORT_mask) begin
      dataArray_3_11[dataArray_3_11_MPORT_addr] <= dataArray_3_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_12_MPORT_en & dataArray_3_12_MPORT_mask) begin
      dataArray_3_12[dataArray_3_12_MPORT_addr] <= dataArray_3_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_13_MPORT_en & dataArray_3_13_MPORT_mask) begin
      dataArray_3_13[dataArray_3_13_MPORT_addr] <= dataArray_3_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_14_MPORT_en & dataArray_3_14_MPORT_mask) begin
      dataArray_3_14[dataArray_3_14_MPORT_addr] <= dataArray_3_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_3_15_MPORT_en & dataArray_3_15_MPORT_mask) begin
      dataArray_3_15[dataArray_3_15_MPORT_addr] <= dataArray_3_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_3_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_3_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_3_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_0_MPORT_en & dataArray_4_0_MPORT_mask) begin
      dataArray_4_0[dataArray_4_0_MPORT_addr] <= dataArray_4_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_1_MPORT_en & dataArray_4_1_MPORT_mask) begin
      dataArray_4_1[dataArray_4_1_MPORT_addr] <= dataArray_4_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_2_MPORT_en & dataArray_4_2_MPORT_mask) begin
      dataArray_4_2[dataArray_4_2_MPORT_addr] <= dataArray_4_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_3_MPORT_en & dataArray_4_3_MPORT_mask) begin
      dataArray_4_3[dataArray_4_3_MPORT_addr] <= dataArray_4_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_4_MPORT_en & dataArray_4_4_MPORT_mask) begin
      dataArray_4_4[dataArray_4_4_MPORT_addr] <= dataArray_4_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_5_MPORT_en & dataArray_4_5_MPORT_mask) begin
      dataArray_4_5[dataArray_4_5_MPORT_addr] <= dataArray_4_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_6_MPORT_en & dataArray_4_6_MPORT_mask) begin
      dataArray_4_6[dataArray_4_6_MPORT_addr] <= dataArray_4_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_7_MPORT_en & dataArray_4_7_MPORT_mask) begin
      dataArray_4_7[dataArray_4_7_MPORT_addr] <= dataArray_4_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_8_MPORT_en & dataArray_4_8_MPORT_mask) begin
      dataArray_4_8[dataArray_4_8_MPORT_addr] <= dataArray_4_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_9_MPORT_en & dataArray_4_9_MPORT_mask) begin
      dataArray_4_9[dataArray_4_9_MPORT_addr] <= dataArray_4_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_10_MPORT_en & dataArray_4_10_MPORT_mask) begin
      dataArray_4_10[dataArray_4_10_MPORT_addr] <= dataArray_4_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_11_MPORT_en & dataArray_4_11_MPORT_mask) begin
      dataArray_4_11[dataArray_4_11_MPORT_addr] <= dataArray_4_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_12_MPORT_en & dataArray_4_12_MPORT_mask) begin
      dataArray_4_12[dataArray_4_12_MPORT_addr] <= dataArray_4_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_13_MPORT_en & dataArray_4_13_MPORT_mask) begin
      dataArray_4_13[dataArray_4_13_MPORT_addr] <= dataArray_4_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_14_MPORT_en & dataArray_4_14_MPORT_mask) begin
      dataArray_4_14[dataArray_4_14_MPORT_addr] <= dataArray_4_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_4_15_MPORT_en & dataArray_4_15_MPORT_mask) begin
      dataArray_4_15[dataArray_4_15_MPORT_addr] <= dataArray_4_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_4_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_4_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_4_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_0_MPORT_en & dataArray_5_0_MPORT_mask) begin
      dataArray_5_0[dataArray_5_0_MPORT_addr] <= dataArray_5_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_1_MPORT_en & dataArray_5_1_MPORT_mask) begin
      dataArray_5_1[dataArray_5_1_MPORT_addr] <= dataArray_5_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_2_MPORT_en & dataArray_5_2_MPORT_mask) begin
      dataArray_5_2[dataArray_5_2_MPORT_addr] <= dataArray_5_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_3_MPORT_en & dataArray_5_3_MPORT_mask) begin
      dataArray_5_3[dataArray_5_3_MPORT_addr] <= dataArray_5_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_4_MPORT_en & dataArray_5_4_MPORT_mask) begin
      dataArray_5_4[dataArray_5_4_MPORT_addr] <= dataArray_5_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_5_MPORT_en & dataArray_5_5_MPORT_mask) begin
      dataArray_5_5[dataArray_5_5_MPORT_addr] <= dataArray_5_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_6_MPORT_en & dataArray_5_6_MPORT_mask) begin
      dataArray_5_6[dataArray_5_6_MPORT_addr] <= dataArray_5_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_7_MPORT_en & dataArray_5_7_MPORT_mask) begin
      dataArray_5_7[dataArray_5_7_MPORT_addr] <= dataArray_5_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_8_MPORT_en & dataArray_5_8_MPORT_mask) begin
      dataArray_5_8[dataArray_5_8_MPORT_addr] <= dataArray_5_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_9_MPORT_en & dataArray_5_9_MPORT_mask) begin
      dataArray_5_9[dataArray_5_9_MPORT_addr] <= dataArray_5_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_10_MPORT_en & dataArray_5_10_MPORT_mask) begin
      dataArray_5_10[dataArray_5_10_MPORT_addr] <= dataArray_5_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_11_MPORT_en & dataArray_5_11_MPORT_mask) begin
      dataArray_5_11[dataArray_5_11_MPORT_addr] <= dataArray_5_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_12_MPORT_en & dataArray_5_12_MPORT_mask) begin
      dataArray_5_12[dataArray_5_12_MPORT_addr] <= dataArray_5_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_13_MPORT_en & dataArray_5_13_MPORT_mask) begin
      dataArray_5_13[dataArray_5_13_MPORT_addr] <= dataArray_5_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_14_MPORT_en & dataArray_5_14_MPORT_mask) begin
      dataArray_5_14[dataArray_5_14_MPORT_addr] <= dataArray_5_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_5_15_MPORT_en & dataArray_5_15_MPORT_mask) begin
      dataArray_5_15[dataArray_5_15_MPORT_addr] <= dataArray_5_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_5_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_5_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_5_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_0_MPORT_en & dataArray_6_0_MPORT_mask) begin
      dataArray_6_0[dataArray_6_0_MPORT_addr] <= dataArray_6_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_1_MPORT_en & dataArray_6_1_MPORT_mask) begin
      dataArray_6_1[dataArray_6_1_MPORT_addr] <= dataArray_6_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_2_MPORT_en & dataArray_6_2_MPORT_mask) begin
      dataArray_6_2[dataArray_6_2_MPORT_addr] <= dataArray_6_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_3_MPORT_en & dataArray_6_3_MPORT_mask) begin
      dataArray_6_3[dataArray_6_3_MPORT_addr] <= dataArray_6_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_4_MPORT_en & dataArray_6_4_MPORT_mask) begin
      dataArray_6_4[dataArray_6_4_MPORT_addr] <= dataArray_6_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_5_MPORT_en & dataArray_6_5_MPORT_mask) begin
      dataArray_6_5[dataArray_6_5_MPORT_addr] <= dataArray_6_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_6_MPORT_en & dataArray_6_6_MPORT_mask) begin
      dataArray_6_6[dataArray_6_6_MPORT_addr] <= dataArray_6_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_7_MPORT_en & dataArray_6_7_MPORT_mask) begin
      dataArray_6_7[dataArray_6_7_MPORT_addr] <= dataArray_6_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_8_MPORT_en & dataArray_6_8_MPORT_mask) begin
      dataArray_6_8[dataArray_6_8_MPORT_addr] <= dataArray_6_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_9_MPORT_en & dataArray_6_9_MPORT_mask) begin
      dataArray_6_9[dataArray_6_9_MPORT_addr] <= dataArray_6_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_10_MPORT_en & dataArray_6_10_MPORT_mask) begin
      dataArray_6_10[dataArray_6_10_MPORT_addr] <= dataArray_6_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_11_MPORT_en & dataArray_6_11_MPORT_mask) begin
      dataArray_6_11[dataArray_6_11_MPORT_addr] <= dataArray_6_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_12_MPORT_en & dataArray_6_12_MPORT_mask) begin
      dataArray_6_12[dataArray_6_12_MPORT_addr] <= dataArray_6_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_13_MPORT_en & dataArray_6_13_MPORT_mask) begin
      dataArray_6_13[dataArray_6_13_MPORT_addr] <= dataArray_6_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_14_MPORT_en & dataArray_6_14_MPORT_mask) begin
      dataArray_6_14[dataArray_6_14_MPORT_addr] <= dataArray_6_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_6_15_MPORT_en & dataArray_6_15_MPORT_mask) begin
      dataArray_6_15[dataArray_6_15_MPORT_addr] <= dataArray_6_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_6_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_6_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_6_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_0_MPORT_en & dataArray_7_0_MPORT_mask) begin
      dataArray_7_0[dataArray_7_0_MPORT_addr] <= dataArray_7_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_1_MPORT_en & dataArray_7_1_MPORT_mask) begin
      dataArray_7_1[dataArray_7_1_MPORT_addr] <= dataArray_7_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_2_MPORT_en & dataArray_7_2_MPORT_mask) begin
      dataArray_7_2[dataArray_7_2_MPORT_addr] <= dataArray_7_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_3_MPORT_en & dataArray_7_3_MPORT_mask) begin
      dataArray_7_3[dataArray_7_3_MPORT_addr] <= dataArray_7_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_4_MPORT_en & dataArray_7_4_MPORT_mask) begin
      dataArray_7_4[dataArray_7_4_MPORT_addr] <= dataArray_7_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_5_MPORT_en & dataArray_7_5_MPORT_mask) begin
      dataArray_7_5[dataArray_7_5_MPORT_addr] <= dataArray_7_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_6_MPORT_en & dataArray_7_6_MPORT_mask) begin
      dataArray_7_6[dataArray_7_6_MPORT_addr] <= dataArray_7_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_7_MPORT_en & dataArray_7_7_MPORT_mask) begin
      dataArray_7_7[dataArray_7_7_MPORT_addr] <= dataArray_7_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_8_MPORT_en & dataArray_7_8_MPORT_mask) begin
      dataArray_7_8[dataArray_7_8_MPORT_addr] <= dataArray_7_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_9_MPORT_en & dataArray_7_9_MPORT_mask) begin
      dataArray_7_9[dataArray_7_9_MPORT_addr] <= dataArray_7_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_10_MPORT_en & dataArray_7_10_MPORT_mask) begin
      dataArray_7_10[dataArray_7_10_MPORT_addr] <= dataArray_7_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_11_MPORT_en & dataArray_7_11_MPORT_mask) begin
      dataArray_7_11[dataArray_7_11_MPORT_addr] <= dataArray_7_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_12_MPORT_en & dataArray_7_12_MPORT_mask) begin
      dataArray_7_12[dataArray_7_12_MPORT_addr] <= dataArray_7_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_13_MPORT_en & dataArray_7_13_MPORT_mask) begin
      dataArray_7_13[dataArray_7_13_MPORT_addr] <= dataArray_7_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_14_MPORT_en & dataArray_7_14_MPORT_mask) begin
      dataArray_7_14[dataArray_7_14_MPORT_addr] <= dataArray_7_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_7_15_MPORT_en & dataArray_7_15_MPORT_mask) begin
      dataArray_7_15[dataArray_7_15_MPORT_addr] <= dataArray_7_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_7_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_7_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_7_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_0_MPORT_en & dataArray_8_0_MPORT_mask) begin
      dataArray_8_0[dataArray_8_0_MPORT_addr] <= dataArray_8_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_1_MPORT_en & dataArray_8_1_MPORT_mask) begin
      dataArray_8_1[dataArray_8_1_MPORT_addr] <= dataArray_8_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_2_MPORT_en & dataArray_8_2_MPORT_mask) begin
      dataArray_8_2[dataArray_8_2_MPORT_addr] <= dataArray_8_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_3_MPORT_en & dataArray_8_3_MPORT_mask) begin
      dataArray_8_3[dataArray_8_3_MPORT_addr] <= dataArray_8_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_4_MPORT_en & dataArray_8_4_MPORT_mask) begin
      dataArray_8_4[dataArray_8_4_MPORT_addr] <= dataArray_8_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_5_MPORT_en & dataArray_8_5_MPORT_mask) begin
      dataArray_8_5[dataArray_8_5_MPORT_addr] <= dataArray_8_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_6_MPORT_en & dataArray_8_6_MPORT_mask) begin
      dataArray_8_6[dataArray_8_6_MPORT_addr] <= dataArray_8_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_7_MPORT_en & dataArray_8_7_MPORT_mask) begin
      dataArray_8_7[dataArray_8_7_MPORT_addr] <= dataArray_8_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_8_MPORT_en & dataArray_8_8_MPORT_mask) begin
      dataArray_8_8[dataArray_8_8_MPORT_addr] <= dataArray_8_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_9_MPORT_en & dataArray_8_9_MPORT_mask) begin
      dataArray_8_9[dataArray_8_9_MPORT_addr] <= dataArray_8_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_10_MPORT_en & dataArray_8_10_MPORT_mask) begin
      dataArray_8_10[dataArray_8_10_MPORT_addr] <= dataArray_8_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_11_MPORT_en & dataArray_8_11_MPORT_mask) begin
      dataArray_8_11[dataArray_8_11_MPORT_addr] <= dataArray_8_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_12_MPORT_en & dataArray_8_12_MPORT_mask) begin
      dataArray_8_12[dataArray_8_12_MPORT_addr] <= dataArray_8_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_13_MPORT_en & dataArray_8_13_MPORT_mask) begin
      dataArray_8_13[dataArray_8_13_MPORT_addr] <= dataArray_8_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_14_MPORT_en & dataArray_8_14_MPORT_mask) begin
      dataArray_8_14[dataArray_8_14_MPORT_addr] <= dataArray_8_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_8_15_MPORT_en & dataArray_8_15_MPORT_mask) begin
      dataArray_8_15[dataArray_8_15_MPORT_addr] <= dataArray_8_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_8_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_8_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_8_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_0_MPORT_en & dataArray_9_0_MPORT_mask) begin
      dataArray_9_0[dataArray_9_0_MPORT_addr] <= dataArray_9_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_1_MPORT_en & dataArray_9_1_MPORT_mask) begin
      dataArray_9_1[dataArray_9_1_MPORT_addr] <= dataArray_9_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_2_MPORT_en & dataArray_9_2_MPORT_mask) begin
      dataArray_9_2[dataArray_9_2_MPORT_addr] <= dataArray_9_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_3_MPORT_en & dataArray_9_3_MPORT_mask) begin
      dataArray_9_3[dataArray_9_3_MPORT_addr] <= dataArray_9_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_4_MPORT_en & dataArray_9_4_MPORT_mask) begin
      dataArray_9_4[dataArray_9_4_MPORT_addr] <= dataArray_9_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_5_MPORT_en & dataArray_9_5_MPORT_mask) begin
      dataArray_9_5[dataArray_9_5_MPORT_addr] <= dataArray_9_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_6_MPORT_en & dataArray_9_6_MPORT_mask) begin
      dataArray_9_6[dataArray_9_6_MPORT_addr] <= dataArray_9_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_7_MPORT_en & dataArray_9_7_MPORT_mask) begin
      dataArray_9_7[dataArray_9_7_MPORT_addr] <= dataArray_9_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_8_MPORT_en & dataArray_9_8_MPORT_mask) begin
      dataArray_9_8[dataArray_9_8_MPORT_addr] <= dataArray_9_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_9_MPORT_en & dataArray_9_9_MPORT_mask) begin
      dataArray_9_9[dataArray_9_9_MPORT_addr] <= dataArray_9_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_10_MPORT_en & dataArray_9_10_MPORT_mask) begin
      dataArray_9_10[dataArray_9_10_MPORT_addr] <= dataArray_9_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_11_MPORT_en & dataArray_9_11_MPORT_mask) begin
      dataArray_9_11[dataArray_9_11_MPORT_addr] <= dataArray_9_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_12_MPORT_en & dataArray_9_12_MPORT_mask) begin
      dataArray_9_12[dataArray_9_12_MPORT_addr] <= dataArray_9_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_13_MPORT_en & dataArray_9_13_MPORT_mask) begin
      dataArray_9_13[dataArray_9_13_MPORT_addr] <= dataArray_9_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_14_MPORT_en & dataArray_9_14_MPORT_mask) begin
      dataArray_9_14[dataArray_9_14_MPORT_addr] <= dataArray_9_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_9_15_MPORT_en & dataArray_9_15_MPORT_mask) begin
      dataArray_9_15[dataArray_9_15_MPORT_addr] <= dataArray_9_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_9_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_9_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_9_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_0_MPORT_en & dataArray_10_0_MPORT_mask) begin
      dataArray_10_0[dataArray_10_0_MPORT_addr] <= dataArray_10_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_1_MPORT_en & dataArray_10_1_MPORT_mask) begin
      dataArray_10_1[dataArray_10_1_MPORT_addr] <= dataArray_10_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_2_MPORT_en & dataArray_10_2_MPORT_mask) begin
      dataArray_10_2[dataArray_10_2_MPORT_addr] <= dataArray_10_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_3_MPORT_en & dataArray_10_3_MPORT_mask) begin
      dataArray_10_3[dataArray_10_3_MPORT_addr] <= dataArray_10_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_4_MPORT_en & dataArray_10_4_MPORT_mask) begin
      dataArray_10_4[dataArray_10_4_MPORT_addr] <= dataArray_10_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_5_MPORT_en & dataArray_10_5_MPORT_mask) begin
      dataArray_10_5[dataArray_10_5_MPORT_addr] <= dataArray_10_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_6_MPORT_en & dataArray_10_6_MPORT_mask) begin
      dataArray_10_6[dataArray_10_6_MPORT_addr] <= dataArray_10_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_7_MPORT_en & dataArray_10_7_MPORT_mask) begin
      dataArray_10_7[dataArray_10_7_MPORT_addr] <= dataArray_10_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_8_MPORT_en & dataArray_10_8_MPORT_mask) begin
      dataArray_10_8[dataArray_10_8_MPORT_addr] <= dataArray_10_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_9_MPORT_en & dataArray_10_9_MPORT_mask) begin
      dataArray_10_9[dataArray_10_9_MPORT_addr] <= dataArray_10_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_10_MPORT_en & dataArray_10_10_MPORT_mask) begin
      dataArray_10_10[dataArray_10_10_MPORT_addr] <= dataArray_10_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_11_MPORT_en & dataArray_10_11_MPORT_mask) begin
      dataArray_10_11[dataArray_10_11_MPORT_addr] <= dataArray_10_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_12_MPORT_en & dataArray_10_12_MPORT_mask) begin
      dataArray_10_12[dataArray_10_12_MPORT_addr] <= dataArray_10_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_13_MPORT_en & dataArray_10_13_MPORT_mask) begin
      dataArray_10_13[dataArray_10_13_MPORT_addr] <= dataArray_10_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_14_MPORT_en & dataArray_10_14_MPORT_mask) begin
      dataArray_10_14[dataArray_10_14_MPORT_addr] <= dataArray_10_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_10_15_MPORT_en & dataArray_10_15_MPORT_mask) begin
      dataArray_10_15[dataArray_10_15_MPORT_addr] <= dataArray_10_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_10_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_10_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_10_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_0_MPORT_en & dataArray_11_0_MPORT_mask) begin
      dataArray_11_0[dataArray_11_0_MPORT_addr] <= dataArray_11_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_1_MPORT_en & dataArray_11_1_MPORT_mask) begin
      dataArray_11_1[dataArray_11_1_MPORT_addr] <= dataArray_11_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_2_MPORT_en & dataArray_11_2_MPORT_mask) begin
      dataArray_11_2[dataArray_11_2_MPORT_addr] <= dataArray_11_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_3_MPORT_en & dataArray_11_3_MPORT_mask) begin
      dataArray_11_3[dataArray_11_3_MPORT_addr] <= dataArray_11_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_4_MPORT_en & dataArray_11_4_MPORT_mask) begin
      dataArray_11_4[dataArray_11_4_MPORT_addr] <= dataArray_11_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_5_MPORT_en & dataArray_11_5_MPORT_mask) begin
      dataArray_11_5[dataArray_11_5_MPORT_addr] <= dataArray_11_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_6_MPORT_en & dataArray_11_6_MPORT_mask) begin
      dataArray_11_6[dataArray_11_6_MPORT_addr] <= dataArray_11_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_7_MPORT_en & dataArray_11_7_MPORT_mask) begin
      dataArray_11_7[dataArray_11_7_MPORT_addr] <= dataArray_11_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_8_MPORT_en & dataArray_11_8_MPORT_mask) begin
      dataArray_11_8[dataArray_11_8_MPORT_addr] <= dataArray_11_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_9_MPORT_en & dataArray_11_9_MPORT_mask) begin
      dataArray_11_9[dataArray_11_9_MPORT_addr] <= dataArray_11_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_10_MPORT_en & dataArray_11_10_MPORT_mask) begin
      dataArray_11_10[dataArray_11_10_MPORT_addr] <= dataArray_11_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_11_MPORT_en & dataArray_11_11_MPORT_mask) begin
      dataArray_11_11[dataArray_11_11_MPORT_addr] <= dataArray_11_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_12_MPORT_en & dataArray_11_12_MPORT_mask) begin
      dataArray_11_12[dataArray_11_12_MPORT_addr] <= dataArray_11_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_13_MPORT_en & dataArray_11_13_MPORT_mask) begin
      dataArray_11_13[dataArray_11_13_MPORT_addr] <= dataArray_11_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_14_MPORT_en & dataArray_11_14_MPORT_mask) begin
      dataArray_11_14[dataArray_11_14_MPORT_addr] <= dataArray_11_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_11_15_MPORT_en & dataArray_11_15_MPORT_mask) begin
      dataArray_11_15[dataArray_11_15_MPORT_addr] <= dataArray_11_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_11_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_11_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_11_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_0_MPORT_en & dataArray_12_0_MPORT_mask) begin
      dataArray_12_0[dataArray_12_0_MPORT_addr] <= dataArray_12_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_1_MPORT_en & dataArray_12_1_MPORT_mask) begin
      dataArray_12_1[dataArray_12_1_MPORT_addr] <= dataArray_12_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_2_MPORT_en & dataArray_12_2_MPORT_mask) begin
      dataArray_12_2[dataArray_12_2_MPORT_addr] <= dataArray_12_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_3_MPORT_en & dataArray_12_3_MPORT_mask) begin
      dataArray_12_3[dataArray_12_3_MPORT_addr] <= dataArray_12_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_4_MPORT_en & dataArray_12_4_MPORT_mask) begin
      dataArray_12_4[dataArray_12_4_MPORT_addr] <= dataArray_12_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_5_MPORT_en & dataArray_12_5_MPORT_mask) begin
      dataArray_12_5[dataArray_12_5_MPORT_addr] <= dataArray_12_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_6_MPORT_en & dataArray_12_6_MPORT_mask) begin
      dataArray_12_6[dataArray_12_6_MPORT_addr] <= dataArray_12_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_7_MPORT_en & dataArray_12_7_MPORT_mask) begin
      dataArray_12_7[dataArray_12_7_MPORT_addr] <= dataArray_12_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_8_MPORT_en & dataArray_12_8_MPORT_mask) begin
      dataArray_12_8[dataArray_12_8_MPORT_addr] <= dataArray_12_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_9_MPORT_en & dataArray_12_9_MPORT_mask) begin
      dataArray_12_9[dataArray_12_9_MPORT_addr] <= dataArray_12_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_10_MPORT_en & dataArray_12_10_MPORT_mask) begin
      dataArray_12_10[dataArray_12_10_MPORT_addr] <= dataArray_12_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_11_MPORT_en & dataArray_12_11_MPORT_mask) begin
      dataArray_12_11[dataArray_12_11_MPORT_addr] <= dataArray_12_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_12_MPORT_en & dataArray_12_12_MPORT_mask) begin
      dataArray_12_12[dataArray_12_12_MPORT_addr] <= dataArray_12_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_13_MPORT_en & dataArray_12_13_MPORT_mask) begin
      dataArray_12_13[dataArray_12_13_MPORT_addr] <= dataArray_12_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_14_MPORT_en & dataArray_12_14_MPORT_mask) begin
      dataArray_12_14[dataArray_12_14_MPORT_addr] <= dataArray_12_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_12_15_MPORT_en & dataArray_12_15_MPORT_mask) begin
      dataArray_12_15[dataArray_12_15_MPORT_addr] <= dataArray_12_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_12_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_12_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_12_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_0_MPORT_en & dataArray_13_0_MPORT_mask) begin
      dataArray_13_0[dataArray_13_0_MPORT_addr] <= dataArray_13_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_1_MPORT_en & dataArray_13_1_MPORT_mask) begin
      dataArray_13_1[dataArray_13_1_MPORT_addr] <= dataArray_13_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_2_MPORT_en & dataArray_13_2_MPORT_mask) begin
      dataArray_13_2[dataArray_13_2_MPORT_addr] <= dataArray_13_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_3_MPORT_en & dataArray_13_3_MPORT_mask) begin
      dataArray_13_3[dataArray_13_3_MPORT_addr] <= dataArray_13_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_4_MPORT_en & dataArray_13_4_MPORT_mask) begin
      dataArray_13_4[dataArray_13_4_MPORT_addr] <= dataArray_13_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_5_MPORT_en & dataArray_13_5_MPORT_mask) begin
      dataArray_13_5[dataArray_13_5_MPORT_addr] <= dataArray_13_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_6_MPORT_en & dataArray_13_6_MPORT_mask) begin
      dataArray_13_6[dataArray_13_6_MPORT_addr] <= dataArray_13_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_7_MPORT_en & dataArray_13_7_MPORT_mask) begin
      dataArray_13_7[dataArray_13_7_MPORT_addr] <= dataArray_13_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_8_MPORT_en & dataArray_13_8_MPORT_mask) begin
      dataArray_13_8[dataArray_13_8_MPORT_addr] <= dataArray_13_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_9_MPORT_en & dataArray_13_9_MPORT_mask) begin
      dataArray_13_9[dataArray_13_9_MPORT_addr] <= dataArray_13_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_10_MPORT_en & dataArray_13_10_MPORT_mask) begin
      dataArray_13_10[dataArray_13_10_MPORT_addr] <= dataArray_13_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_11_MPORT_en & dataArray_13_11_MPORT_mask) begin
      dataArray_13_11[dataArray_13_11_MPORT_addr] <= dataArray_13_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_12_MPORT_en & dataArray_13_12_MPORT_mask) begin
      dataArray_13_12[dataArray_13_12_MPORT_addr] <= dataArray_13_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_13_MPORT_en & dataArray_13_13_MPORT_mask) begin
      dataArray_13_13[dataArray_13_13_MPORT_addr] <= dataArray_13_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_14_MPORT_en & dataArray_13_14_MPORT_mask) begin
      dataArray_13_14[dataArray_13_14_MPORT_addr] <= dataArray_13_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_13_15_MPORT_en & dataArray_13_15_MPORT_mask) begin
      dataArray_13_15[dataArray_13_15_MPORT_addr] <= dataArray_13_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_13_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_13_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_13_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_0_MPORT_en & dataArray_14_0_MPORT_mask) begin
      dataArray_14_0[dataArray_14_0_MPORT_addr] <= dataArray_14_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_1_MPORT_en & dataArray_14_1_MPORT_mask) begin
      dataArray_14_1[dataArray_14_1_MPORT_addr] <= dataArray_14_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_2_MPORT_en & dataArray_14_2_MPORT_mask) begin
      dataArray_14_2[dataArray_14_2_MPORT_addr] <= dataArray_14_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_3_MPORT_en & dataArray_14_3_MPORT_mask) begin
      dataArray_14_3[dataArray_14_3_MPORT_addr] <= dataArray_14_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_4_MPORT_en & dataArray_14_4_MPORT_mask) begin
      dataArray_14_4[dataArray_14_4_MPORT_addr] <= dataArray_14_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_5_MPORT_en & dataArray_14_5_MPORT_mask) begin
      dataArray_14_5[dataArray_14_5_MPORT_addr] <= dataArray_14_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_6_MPORT_en & dataArray_14_6_MPORT_mask) begin
      dataArray_14_6[dataArray_14_6_MPORT_addr] <= dataArray_14_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_7_MPORT_en & dataArray_14_7_MPORT_mask) begin
      dataArray_14_7[dataArray_14_7_MPORT_addr] <= dataArray_14_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_8_MPORT_en & dataArray_14_8_MPORT_mask) begin
      dataArray_14_8[dataArray_14_8_MPORT_addr] <= dataArray_14_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_9_MPORT_en & dataArray_14_9_MPORT_mask) begin
      dataArray_14_9[dataArray_14_9_MPORT_addr] <= dataArray_14_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_10_MPORT_en & dataArray_14_10_MPORT_mask) begin
      dataArray_14_10[dataArray_14_10_MPORT_addr] <= dataArray_14_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_11_MPORT_en & dataArray_14_11_MPORT_mask) begin
      dataArray_14_11[dataArray_14_11_MPORT_addr] <= dataArray_14_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_12_MPORT_en & dataArray_14_12_MPORT_mask) begin
      dataArray_14_12[dataArray_14_12_MPORT_addr] <= dataArray_14_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_13_MPORT_en & dataArray_14_13_MPORT_mask) begin
      dataArray_14_13[dataArray_14_13_MPORT_addr] <= dataArray_14_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_14_MPORT_en & dataArray_14_14_MPORT_mask) begin
      dataArray_14_14[dataArray_14_14_MPORT_addr] <= dataArray_14_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_14_15_MPORT_en & dataArray_14_15_MPORT_mask) begin
      dataArray_14_15[dataArray_14_15_MPORT_addr] <= dataArray_14_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_14_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_14_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_14_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_0_MPORT_en & dataArray_15_0_MPORT_mask) begin
      dataArray_15_0[dataArray_15_0_MPORT_addr] <= dataArray_15_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_1_MPORT_en & dataArray_15_1_MPORT_mask) begin
      dataArray_15_1[dataArray_15_1_MPORT_addr] <= dataArray_15_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_2_MPORT_en & dataArray_15_2_MPORT_mask) begin
      dataArray_15_2[dataArray_15_2_MPORT_addr] <= dataArray_15_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_3_MPORT_en & dataArray_15_3_MPORT_mask) begin
      dataArray_15_3[dataArray_15_3_MPORT_addr] <= dataArray_15_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_4_MPORT_en & dataArray_15_4_MPORT_mask) begin
      dataArray_15_4[dataArray_15_4_MPORT_addr] <= dataArray_15_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_5_MPORT_en & dataArray_15_5_MPORT_mask) begin
      dataArray_15_5[dataArray_15_5_MPORT_addr] <= dataArray_15_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_6_MPORT_en & dataArray_15_6_MPORT_mask) begin
      dataArray_15_6[dataArray_15_6_MPORT_addr] <= dataArray_15_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_7_MPORT_en & dataArray_15_7_MPORT_mask) begin
      dataArray_15_7[dataArray_15_7_MPORT_addr] <= dataArray_15_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_8_MPORT_en & dataArray_15_8_MPORT_mask) begin
      dataArray_15_8[dataArray_15_8_MPORT_addr] <= dataArray_15_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_9_MPORT_en & dataArray_15_9_MPORT_mask) begin
      dataArray_15_9[dataArray_15_9_MPORT_addr] <= dataArray_15_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_10_MPORT_en & dataArray_15_10_MPORT_mask) begin
      dataArray_15_10[dataArray_15_10_MPORT_addr] <= dataArray_15_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_11_MPORT_en & dataArray_15_11_MPORT_mask) begin
      dataArray_15_11[dataArray_15_11_MPORT_addr] <= dataArray_15_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_12_MPORT_en & dataArray_15_12_MPORT_mask) begin
      dataArray_15_12[dataArray_15_12_MPORT_addr] <= dataArray_15_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_13_MPORT_en & dataArray_15_13_MPORT_mask) begin
      dataArray_15_13[dataArray_15_13_MPORT_addr] <= dataArray_15_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_14_MPORT_en & dataArray_15_14_MPORT_mask) begin
      dataArray_15_14[dataArray_15_14_MPORT_addr] <= dataArray_15_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_15_15_MPORT_en & dataArray_15_15_MPORT_mask) begin
      dataArray_15_15[dataArray_15_15_MPORT_addr] <= dataArray_15_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_15_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_15_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_15_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_0_MPORT_en & dataArray_16_0_MPORT_mask) begin
      dataArray_16_0[dataArray_16_0_MPORT_addr] <= dataArray_16_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_1_MPORT_en & dataArray_16_1_MPORT_mask) begin
      dataArray_16_1[dataArray_16_1_MPORT_addr] <= dataArray_16_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_2_MPORT_en & dataArray_16_2_MPORT_mask) begin
      dataArray_16_2[dataArray_16_2_MPORT_addr] <= dataArray_16_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_3_MPORT_en & dataArray_16_3_MPORT_mask) begin
      dataArray_16_3[dataArray_16_3_MPORT_addr] <= dataArray_16_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_4_MPORT_en & dataArray_16_4_MPORT_mask) begin
      dataArray_16_4[dataArray_16_4_MPORT_addr] <= dataArray_16_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_5_MPORT_en & dataArray_16_5_MPORT_mask) begin
      dataArray_16_5[dataArray_16_5_MPORT_addr] <= dataArray_16_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_6_MPORT_en & dataArray_16_6_MPORT_mask) begin
      dataArray_16_6[dataArray_16_6_MPORT_addr] <= dataArray_16_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_7_MPORT_en & dataArray_16_7_MPORT_mask) begin
      dataArray_16_7[dataArray_16_7_MPORT_addr] <= dataArray_16_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_8_MPORT_en & dataArray_16_8_MPORT_mask) begin
      dataArray_16_8[dataArray_16_8_MPORT_addr] <= dataArray_16_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_9_MPORT_en & dataArray_16_9_MPORT_mask) begin
      dataArray_16_9[dataArray_16_9_MPORT_addr] <= dataArray_16_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_10_MPORT_en & dataArray_16_10_MPORT_mask) begin
      dataArray_16_10[dataArray_16_10_MPORT_addr] <= dataArray_16_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_11_MPORT_en & dataArray_16_11_MPORT_mask) begin
      dataArray_16_11[dataArray_16_11_MPORT_addr] <= dataArray_16_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_12_MPORT_en & dataArray_16_12_MPORT_mask) begin
      dataArray_16_12[dataArray_16_12_MPORT_addr] <= dataArray_16_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_13_MPORT_en & dataArray_16_13_MPORT_mask) begin
      dataArray_16_13[dataArray_16_13_MPORT_addr] <= dataArray_16_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_14_MPORT_en & dataArray_16_14_MPORT_mask) begin
      dataArray_16_14[dataArray_16_14_MPORT_addr] <= dataArray_16_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_16_15_MPORT_en & dataArray_16_15_MPORT_mask) begin
      dataArray_16_15[dataArray_16_15_MPORT_addr] <= dataArray_16_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_16_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_16_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_16_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_16_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_0_MPORT_en & dataArray_17_0_MPORT_mask) begin
      dataArray_17_0[dataArray_17_0_MPORT_addr] <= dataArray_17_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_1_MPORT_en & dataArray_17_1_MPORT_mask) begin
      dataArray_17_1[dataArray_17_1_MPORT_addr] <= dataArray_17_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_2_MPORT_en & dataArray_17_2_MPORT_mask) begin
      dataArray_17_2[dataArray_17_2_MPORT_addr] <= dataArray_17_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_3_MPORT_en & dataArray_17_3_MPORT_mask) begin
      dataArray_17_3[dataArray_17_3_MPORT_addr] <= dataArray_17_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_4_MPORT_en & dataArray_17_4_MPORT_mask) begin
      dataArray_17_4[dataArray_17_4_MPORT_addr] <= dataArray_17_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_5_MPORT_en & dataArray_17_5_MPORT_mask) begin
      dataArray_17_5[dataArray_17_5_MPORT_addr] <= dataArray_17_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_6_MPORT_en & dataArray_17_6_MPORT_mask) begin
      dataArray_17_6[dataArray_17_6_MPORT_addr] <= dataArray_17_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_7_MPORT_en & dataArray_17_7_MPORT_mask) begin
      dataArray_17_7[dataArray_17_7_MPORT_addr] <= dataArray_17_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_8_MPORT_en & dataArray_17_8_MPORT_mask) begin
      dataArray_17_8[dataArray_17_8_MPORT_addr] <= dataArray_17_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_9_MPORT_en & dataArray_17_9_MPORT_mask) begin
      dataArray_17_9[dataArray_17_9_MPORT_addr] <= dataArray_17_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_10_MPORT_en & dataArray_17_10_MPORT_mask) begin
      dataArray_17_10[dataArray_17_10_MPORT_addr] <= dataArray_17_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_11_MPORT_en & dataArray_17_11_MPORT_mask) begin
      dataArray_17_11[dataArray_17_11_MPORT_addr] <= dataArray_17_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_12_MPORT_en & dataArray_17_12_MPORT_mask) begin
      dataArray_17_12[dataArray_17_12_MPORT_addr] <= dataArray_17_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_13_MPORT_en & dataArray_17_13_MPORT_mask) begin
      dataArray_17_13[dataArray_17_13_MPORT_addr] <= dataArray_17_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_14_MPORT_en & dataArray_17_14_MPORT_mask) begin
      dataArray_17_14[dataArray_17_14_MPORT_addr] <= dataArray_17_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_17_15_MPORT_en & dataArray_17_15_MPORT_mask) begin
      dataArray_17_15[dataArray_17_15_MPORT_addr] <= dataArray_17_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_17_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_17_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_17_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_17_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_0_MPORT_en & dataArray_18_0_MPORT_mask) begin
      dataArray_18_0[dataArray_18_0_MPORT_addr] <= dataArray_18_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_1_MPORT_en & dataArray_18_1_MPORT_mask) begin
      dataArray_18_1[dataArray_18_1_MPORT_addr] <= dataArray_18_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_2_MPORT_en & dataArray_18_2_MPORT_mask) begin
      dataArray_18_2[dataArray_18_2_MPORT_addr] <= dataArray_18_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_3_MPORT_en & dataArray_18_3_MPORT_mask) begin
      dataArray_18_3[dataArray_18_3_MPORT_addr] <= dataArray_18_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_4_MPORT_en & dataArray_18_4_MPORT_mask) begin
      dataArray_18_4[dataArray_18_4_MPORT_addr] <= dataArray_18_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_5_MPORT_en & dataArray_18_5_MPORT_mask) begin
      dataArray_18_5[dataArray_18_5_MPORT_addr] <= dataArray_18_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_6_MPORT_en & dataArray_18_6_MPORT_mask) begin
      dataArray_18_6[dataArray_18_6_MPORT_addr] <= dataArray_18_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_7_MPORT_en & dataArray_18_7_MPORT_mask) begin
      dataArray_18_7[dataArray_18_7_MPORT_addr] <= dataArray_18_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_8_MPORT_en & dataArray_18_8_MPORT_mask) begin
      dataArray_18_8[dataArray_18_8_MPORT_addr] <= dataArray_18_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_9_MPORT_en & dataArray_18_9_MPORT_mask) begin
      dataArray_18_9[dataArray_18_9_MPORT_addr] <= dataArray_18_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_10_MPORT_en & dataArray_18_10_MPORT_mask) begin
      dataArray_18_10[dataArray_18_10_MPORT_addr] <= dataArray_18_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_11_MPORT_en & dataArray_18_11_MPORT_mask) begin
      dataArray_18_11[dataArray_18_11_MPORT_addr] <= dataArray_18_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_12_MPORT_en & dataArray_18_12_MPORT_mask) begin
      dataArray_18_12[dataArray_18_12_MPORT_addr] <= dataArray_18_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_13_MPORT_en & dataArray_18_13_MPORT_mask) begin
      dataArray_18_13[dataArray_18_13_MPORT_addr] <= dataArray_18_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_14_MPORT_en & dataArray_18_14_MPORT_mask) begin
      dataArray_18_14[dataArray_18_14_MPORT_addr] <= dataArray_18_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_18_15_MPORT_en & dataArray_18_15_MPORT_mask) begin
      dataArray_18_15[dataArray_18_15_MPORT_addr] <= dataArray_18_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_18_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_18_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_18_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_18_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_0_MPORT_en & dataArray_19_0_MPORT_mask) begin
      dataArray_19_0[dataArray_19_0_MPORT_addr] <= dataArray_19_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_1_MPORT_en & dataArray_19_1_MPORT_mask) begin
      dataArray_19_1[dataArray_19_1_MPORT_addr] <= dataArray_19_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_2_MPORT_en & dataArray_19_2_MPORT_mask) begin
      dataArray_19_2[dataArray_19_2_MPORT_addr] <= dataArray_19_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_3_MPORT_en & dataArray_19_3_MPORT_mask) begin
      dataArray_19_3[dataArray_19_3_MPORT_addr] <= dataArray_19_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_4_MPORT_en & dataArray_19_4_MPORT_mask) begin
      dataArray_19_4[dataArray_19_4_MPORT_addr] <= dataArray_19_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_5_MPORT_en & dataArray_19_5_MPORT_mask) begin
      dataArray_19_5[dataArray_19_5_MPORT_addr] <= dataArray_19_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_6_MPORT_en & dataArray_19_6_MPORT_mask) begin
      dataArray_19_6[dataArray_19_6_MPORT_addr] <= dataArray_19_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_7_MPORT_en & dataArray_19_7_MPORT_mask) begin
      dataArray_19_7[dataArray_19_7_MPORT_addr] <= dataArray_19_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_8_MPORT_en & dataArray_19_8_MPORT_mask) begin
      dataArray_19_8[dataArray_19_8_MPORT_addr] <= dataArray_19_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_9_MPORT_en & dataArray_19_9_MPORT_mask) begin
      dataArray_19_9[dataArray_19_9_MPORT_addr] <= dataArray_19_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_10_MPORT_en & dataArray_19_10_MPORT_mask) begin
      dataArray_19_10[dataArray_19_10_MPORT_addr] <= dataArray_19_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_11_MPORT_en & dataArray_19_11_MPORT_mask) begin
      dataArray_19_11[dataArray_19_11_MPORT_addr] <= dataArray_19_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_12_MPORT_en & dataArray_19_12_MPORT_mask) begin
      dataArray_19_12[dataArray_19_12_MPORT_addr] <= dataArray_19_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_13_MPORT_en & dataArray_19_13_MPORT_mask) begin
      dataArray_19_13[dataArray_19_13_MPORT_addr] <= dataArray_19_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_14_MPORT_en & dataArray_19_14_MPORT_mask) begin
      dataArray_19_14[dataArray_19_14_MPORT_addr] <= dataArray_19_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_19_15_MPORT_en & dataArray_19_15_MPORT_mask) begin
      dataArray_19_15[dataArray_19_15_MPORT_addr] <= dataArray_19_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_19_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_19_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_19_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_19_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_0_MPORT_en & dataArray_20_0_MPORT_mask) begin
      dataArray_20_0[dataArray_20_0_MPORT_addr] <= dataArray_20_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_1_MPORT_en & dataArray_20_1_MPORT_mask) begin
      dataArray_20_1[dataArray_20_1_MPORT_addr] <= dataArray_20_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_2_MPORT_en & dataArray_20_2_MPORT_mask) begin
      dataArray_20_2[dataArray_20_2_MPORT_addr] <= dataArray_20_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_3_MPORT_en & dataArray_20_3_MPORT_mask) begin
      dataArray_20_3[dataArray_20_3_MPORT_addr] <= dataArray_20_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_4_MPORT_en & dataArray_20_4_MPORT_mask) begin
      dataArray_20_4[dataArray_20_4_MPORT_addr] <= dataArray_20_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_5_MPORT_en & dataArray_20_5_MPORT_mask) begin
      dataArray_20_5[dataArray_20_5_MPORT_addr] <= dataArray_20_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_6_MPORT_en & dataArray_20_6_MPORT_mask) begin
      dataArray_20_6[dataArray_20_6_MPORT_addr] <= dataArray_20_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_7_MPORT_en & dataArray_20_7_MPORT_mask) begin
      dataArray_20_7[dataArray_20_7_MPORT_addr] <= dataArray_20_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_8_MPORT_en & dataArray_20_8_MPORT_mask) begin
      dataArray_20_8[dataArray_20_8_MPORT_addr] <= dataArray_20_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_9_MPORT_en & dataArray_20_9_MPORT_mask) begin
      dataArray_20_9[dataArray_20_9_MPORT_addr] <= dataArray_20_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_10_MPORT_en & dataArray_20_10_MPORT_mask) begin
      dataArray_20_10[dataArray_20_10_MPORT_addr] <= dataArray_20_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_11_MPORT_en & dataArray_20_11_MPORT_mask) begin
      dataArray_20_11[dataArray_20_11_MPORT_addr] <= dataArray_20_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_12_MPORT_en & dataArray_20_12_MPORT_mask) begin
      dataArray_20_12[dataArray_20_12_MPORT_addr] <= dataArray_20_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_13_MPORT_en & dataArray_20_13_MPORT_mask) begin
      dataArray_20_13[dataArray_20_13_MPORT_addr] <= dataArray_20_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_14_MPORT_en & dataArray_20_14_MPORT_mask) begin
      dataArray_20_14[dataArray_20_14_MPORT_addr] <= dataArray_20_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_20_15_MPORT_en & dataArray_20_15_MPORT_mask) begin
      dataArray_20_15[dataArray_20_15_MPORT_addr] <= dataArray_20_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_20_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_20_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_20_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_20_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_0_MPORT_en & dataArray_21_0_MPORT_mask) begin
      dataArray_21_0[dataArray_21_0_MPORT_addr] <= dataArray_21_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_1_MPORT_en & dataArray_21_1_MPORT_mask) begin
      dataArray_21_1[dataArray_21_1_MPORT_addr] <= dataArray_21_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_2_MPORT_en & dataArray_21_2_MPORT_mask) begin
      dataArray_21_2[dataArray_21_2_MPORT_addr] <= dataArray_21_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_3_MPORT_en & dataArray_21_3_MPORT_mask) begin
      dataArray_21_3[dataArray_21_3_MPORT_addr] <= dataArray_21_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_4_MPORT_en & dataArray_21_4_MPORT_mask) begin
      dataArray_21_4[dataArray_21_4_MPORT_addr] <= dataArray_21_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_5_MPORT_en & dataArray_21_5_MPORT_mask) begin
      dataArray_21_5[dataArray_21_5_MPORT_addr] <= dataArray_21_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_6_MPORT_en & dataArray_21_6_MPORT_mask) begin
      dataArray_21_6[dataArray_21_6_MPORT_addr] <= dataArray_21_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_7_MPORT_en & dataArray_21_7_MPORT_mask) begin
      dataArray_21_7[dataArray_21_7_MPORT_addr] <= dataArray_21_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_8_MPORT_en & dataArray_21_8_MPORT_mask) begin
      dataArray_21_8[dataArray_21_8_MPORT_addr] <= dataArray_21_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_9_MPORT_en & dataArray_21_9_MPORT_mask) begin
      dataArray_21_9[dataArray_21_9_MPORT_addr] <= dataArray_21_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_10_MPORT_en & dataArray_21_10_MPORT_mask) begin
      dataArray_21_10[dataArray_21_10_MPORT_addr] <= dataArray_21_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_11_MPORT_en & dataArray_21_11_MPORT_mask) begin
      dataArray_21_11[dataArray_21_11_MPORT_addr] <= dataArray_21_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_12_MPORT_en & dataArray_21_12_MPORT_mask) begin
      dataArray_21_12[dataArray_21_12_MPORT_addr] <= dataArray_21_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_13_MPORT_en & dataArray_21_13_MPORT_mask) begin
      dataArray_21_13[dataArray_21_13_MPORT_addr] <= dataArray_21_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_14_MPORT_en & dataArray_21_14_MPORT_mask) begin
      dataArray_21_14[dataArray_21_14_MPORT_addr] <= dataArray_21_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_21_15_MPORT_en & dataArray_21_15_MPORT_mask) begin
      dataArray_21_15[dataArray_21_15_MPORT_addr] <= dataArray_21_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_21_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_21_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_21_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_21_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_0_MPORT_en & dataArray_22_0_MPORT_mask) begin
      dataArray_22_0[dataArray_22_0_MPORT_addr] <= dataArray_22_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_1_MPORT_en & dataArray_22_1_MPORT_mask) begin
      dataArray_22_1[dataArray_22_1_MPORT_addr] <= dataArray_22_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_2_MPORT_en & dataArray_22_2_MPORT_mask) begin
      dataArray_22_2[dataArray_22_2_MPORT_addr] <= dataArray_22_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_3_MPORT_en & dataArray_22_3_MPORT_mask) begin
      dataArray_22_3[dataArray_22_3_MPORT_addr] <= dataArray_22_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_4_MPORT_en & dataArray_22_4_MPORT_mask) begin
      dataArray_22_4[dataArray_22_4_MPORT_addr] <= dataArray_22_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_5_MPORT_en & dataArray_22_5_MPORT_mask) begin
      dataArray_22_5[dataArray_22_5_MPORT_addr] <= dataArray_22_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_6_MPORT_en & dataArray_22_6_MPORT_mask) begin
      dataArray_22_6[dataArray_22_6_MPORT_addr] <= dataArray_22_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_7_MPORT_en & dataArray_22_7_MPORT_mask) begin
      dataArray_22_7[dataArray_22_7_MPORT_addr] <= dataArray_22_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_8_MPORT_en & dataArray_22_8_MPORT_mask) begin
      dataArray_22_8[dataArray_22_8_MPORT_addr] <= dataArray_22_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_9_MPORT_en & dataArray_22_9_MPORT_mask) begin
      dataArray_22_9[dataArray_22_9_MPORT_addr] <= dataArray_22_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_10_MPORT_en & dataArray_22_10_MPORT_mask) begin
      dataArray_22_10[dataArray_22_10_MPORT_addr] <= dataArray_22_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_11_MPORT_en & dataArray_22_11_MPORT_mask) begin
      dataArray_22_11[dataArray_22_11_MPORT_addr] <= dataArray_22_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_12_MPORT_en & dataArray_22_12_MPORT_mask) begin
      dataArray_22_12[dataArray_22_12_MPORT_addr] <= dataArray_22_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_13_MPORT_en & dataArray_22_13_MPORT_mask) begin
      dataArray_22_13[dataArray_22_13_MPORT_addr] <= dataArray_22_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_14_MPORT_en & dataArray_22_14_MPORT_mask) begin
      dataArray_22_14[dataArray_22_14_MPORT_addr] <= dataArray_22_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_22_15_MPORT_en & dataArray_22_15_MPORT_mask) begin
      dataArray_22_15[dataArray_22_15_MPORT_addr] <= dataArray_22_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_22_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_22_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_22_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_22_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_0_MPORT_en & dataArray_23_0_MPORT_mask) begin
      dataArray_23_0[dataArray_23_0_MPORT_addr] <= dataArray_23_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_1_MPORT_en & dataArray_23_1_MPORT_mask) begin
      dataArray_23_1[dataArray_23_1_MPORT_addr] <= dataArray_23_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_2_MPORT_en & dataArray_23_2_MPORT_mask) begin
      dataArray_23_2[dataArray_23_2_MPORT_addr] <= dataArray_23_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_3_MPORT_en & dataArray_23_3_MPORT_mask) begin
      dataArray_23_3[dataArray_23_3_MPORT_addr] <= dataArray_23_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_4_MPORT_en & dataArray_23_4_MPORT_mask) begin
      dataArray_23_4[dataArray_23_4_MPORT_addr] <= dataArray_23_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_5_MPORT_en & dataArray_23_5_MPORT_mask) begin
      dataArray_23_5[dataArray_23_5_MPORT_addr] <= dataArray_23_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_6_MPORT_en & dataArray_23_6_MPORT_mask) begin
      dataArray_23_6[dataArray_23_6_MPORT_addr] <= dataArray_23_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_7_MPORT_en & dataArray_23_7_MPORT_mask) begin
      dataArray_23_7[dataArray_23_7_MPORT_addr] <= dataArray_23_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_8_MPORT_en & dataArray_23_8_MPORT_mask) begin
      dataArray_23_8[dataArray_23_8_MPORT_addr] <= dataArray_23_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_9_MPORT_en & dataArray_23_9_MPORT_mask) begin
      dataArray_23_9[dataArray_23_9_MPORT_addr] <= dataArray_23_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_10_MPORT_en & dataArray_23_10_MPORT_mask) begin
      dataArray_23_10[dataArray_23_10_MPORT_addr] <= dataArray_23_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_11_MPORT_en & dataArray_23_11_MPORT_mask) begin
      dataArray_23_11[dataArray_23_11_MPORT_addr] <= dataArray_23_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_12_MPORT_en & dataArray_23_12_MPORT_mask) begin
      dataArray_23_12[dataArray_23_12_MPORT_addr] <= dataArray_23_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_13_MPORT_en & dataArray_23_13_MPORT_mask) begin
      dataArray_23_13[dataArray_23_13_MPORT_addr] <= dataArray_23_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_14_MPORT_en & dataArray_23_14_MPORT_mask) begin
      dataArray_23_14[dataArray_23_14_MPORT_addr] <= dataArray_23_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_23_15_MPORT_en & dataArray_23_15_MPORT_mask) begin
      dataArray_23_15[dataArray_23_15_MPORT_addr] <= dataArray_23_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_23_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_23_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_23_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_23_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_0_MPORT_en & dataArray_24_0_MPORT_mask) begin
      dataArray_24_0[dataArray_24_0_MPORT_addr] <= dataArray_24_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_1_MPORT_en & dataArray_24_1_MPORT_mask) begin
      dataArray_24_1[dataArray_24_1_MPORT_addr] <= dataArray_24_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_2_MPORT_en & dataArray_24_2_MPORT_mask) begin
      dataArray_24_2[dataArray_24_2_MPORT_addr] <= dataArray_24_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_3_MPORT_en & dataArray_24_3_MPORT_mask) begin
      dataArray_24_3[dataArray_24_3_MPORT_addr] <= dataArray_24_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_4_MPORT_en & dataArray_24_4_MPORT_mask) begin
      dataArray_24_4[dataArray_24_4_MPORT_addr] <= dataArray_24_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_5_MPORT_en & dataArray_24_5_MPORT_mask) begin
      dataArray_24_5[dataArray_24_5_MPORT_addr] <= dataArray_24_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_6_MPORT_en & dataArray_24_6_MPORT_mask) begin
      dataArray_24_6[dataArray_24_6_MPORT_addr] <= dataArray_24_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_7_MPORT_en & dataArray_24_7_MPORT_mask) begin
      dataArray_24_7[dataArray_24_7_MPORT_addr] <= dataArray_24_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_8_MPORT_en & dataArray_24_8_MPORT_mask) begin
      dataArray_24_8[dataArray_24_8_MPORT_addr] <= dataArray_24_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_9_MPORT_en & dataArray_24_9_MPORT_mask) begin
      dataArray_24_9[dataArray_24_9_MPORT_addr] <= dataArray_24_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_10_MPORT_en & dataArray_24_10_MPORT_mask) begin
      dataArray_24_10[dataArray_24_10_MPORT_addr] <= dataArray_24_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_11_MPORT_en & dataArray_24_11_MPORT_mask) begin
      dataArray_24_11[dataArray_24_11_MPORT_addr] <= dataArray_24_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_12_MPORT_en & dataArray_24_12_MPORT_mask) begin
      dataArray_24_12[dataArray_24_12_MPORT_addr] <= dataArray_24_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_13_MPORT_en & dataArray_24_13_MPORT_mask) begin
      dataArray_24_13[dataArray_24_13_MPORT_addr] <= dataArray_24_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_14_MPORT_en & dataArray_24_14_MPORT_mask) begin
      dataArray_24_14[dataArray_24_14_MPORT_addr] <= dataArray_24_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_24_15_MPORT_en & dataArray_24_15_MPORT_mask) begin
      dataArray_24_15[dataArray_24_15_MPORT_addr] <= dataArray_24_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_24_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_24_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_24_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_24_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_0_MPORT_en & dataArray_25_0_MPORT_mask) begin
      dataArray_25_0[dataArray_25_0_MPORT_addr] <= dataArray_25_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_1_MPORT_en & dataArray_25_1_MPORT_mask) begin
      dataArray_25_1[dataArray_25_1_MPORT_addr] <= dataArray_25_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_2_MPORT_en & dataArray_25_2_MPORT_mask) begin
      dataArray_25_2[dataArray_25_2_MPORT_addr] <= dataArray_25_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_3_MPORT_en & dataArray_25_3_MPORT_mask) begin
      dataArray_25_3[dataArray_25_3_MPORT_addr] <= dataArray_25_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_4_MPORT_en & dataArray_25_4_MPORT_mask) begin
      dataArray_25_4[dataArray_25_4_MPORT_addr] <= dataArray_25_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_5_MPORT_en & dataArray_25_5_MPORT_mask) begin
      dataArray_25_5[dataArray_25_5_MPORT_addr] <= dataArray_25_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_6_MPORT_en & dataArray_25_6_MPORT_mask) begin
      dataArray_25_6[dataArray_25_6_MPORT_addr] <= dataArray_25_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_7_MPORT_en & dataArray_25_7_MPORT_mask) begin
      dataArray_25_7[dataArray_25_7_MPORT_addr] <= dataArray_25_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_8_MPORT_en & dataArray_25_8_MPORT_mask) begin
      dataArray_25_8[dataArray_25_8_MPORT_addr] <= dataArray_25_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_9_MPORT_en & dataArray_25_9_MPORT_mask) begin
      dataArray_25_9[dataArray_25_9_MPORT_addr] <= dataArray_25_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_10_MPORT_en & dataArray_25_10_MPORT_mask) begin
      dataArray_25_10[dataArray_25_10_MPORT_addr] <= dataArray_25_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_11_MPORT_en & dataArray_25_11_MPORT_mask) begin
      dataArray_25_11[dataArray_25_11_MPORT_addr] <= dataArray_25_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_12_MPORT_en & dataArray_25_12_MPORT_mask) begin
      dataArray_25_12[dataArray_25_12_MPORT_addr] <= dataArray_25_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_13_MPORT_en & dataArray_25_13_MPORT_mask) begin
      dataArray_25_13[dataArray_25_13_MPORT_addr] <= dataArray_25_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_14_MPORT_en & dataArray_25_14_MPORT_mask) begin
      dataArray_25_14[dataArray_25_14_MPORT_addr] <= dataArray_25_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_25_15_MPORT_en & dataArray_25_15_MPORT_mask) begin
      dataArray_25_15[dataArray_25_15_MPORT_addr] <= dataArray_25_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_25_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_25_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_25_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_25_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_0_MPORT_en & dataArray_26_0_MPORT_mask) begin
      dataArray_26_0[dataArray_26_0_MPORT_addr] <= dataArray_26_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_1_MPORT_en & dataArray_26_1_MPORT_mask) begin
      dataArray_26_1[dataArray_26_1_MPORT_addr] <= dataArray_26_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_2_MPORT_en & dataArray_26_2_MPORT_mask) begin
      dataArray_26_2[dataArray_26_2_MPORT_addr] <= dataArray_26_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_3_MPORT_en & dataArray_26_3_MPORT_mask) begin
      dataArray_26_3[dataArray_26_3_MPORT_addr] <= dataArray_26_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_4_MPORT_en & dataArray_26_4_MPORT_mask) begin
      dataArray_26_4[dataArray_26_4_MPORT_addr] <= dataArray_26_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_5_MPORT_en & dataArray_26_5_MPORT_mask) begin
      dataArray_26_5[dataArray_26_5_MPORT_addr] <= dataArray_26_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_6_MPORT_en & dataArray_26_6_MPORT_mask) begin
      dataArray_26_6[dataArray_26_6_MPORT_addr] <= dataArray_26_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_7_MPORT_en & dataArray_26_7_MPORT_mask) begin
      dataArray_26_7[dataArray_26_7_MPORT_addr] <= dataArray_26_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_8_MPORT_en & dataArray_26_8_MPORT_mask) begin
      dataArray_26_8[dataArray_26_8_MPORT_addr] <= dataArray_26_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_9_MPORT_en & dataArray_26_9_MPORT_mask) begin
      dataArray_26_9[dataArray_26_9_MPORT_addr] <= dataArray_26_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_10_MPORT_en & dataArray_26_10_MPORT_mask) begin
      dataArray_26_10[dataArray_26_10_MPORT_addr] <= dataArray_26_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_11_MPORT_en & dataArray_26_11_MPORT_mask) begin
      dataArray_26_11[dataArray_26_11_MPORT_addr] <= dataArray_26_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_12_MPORT_en & dataArray_26_12_MPORT_mask) begin
      dataArray_26_12[dataArray_26_12_MPORT_addr] <= dataArray_26_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_13_MPORT_en & dataArray_26_13_MPORT_mask) begin
      dataArray_26_13[dataArray_26_13_MPORT_addr] <= dataArray_26_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_14_MPORT_en & dataArray_26_14_MPORT_mask) begin
      dataArray_26_14[dataArray_26_14_MPORT_addr] <= dataArray_26_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_26_15_MPORT_en & dataArray_26_15_MPORT_mask) begin
      dataArray_26_15[dataArray_26_15_MPORT_addr] <= dataArray_26_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_26_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_26_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_26_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_26_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_0_MPORT_en & dataArray_27_0_MPORT_mask) begin
      dataArray_27_0[dataArray_27_0_MPORT_addr] <= dataArray_27_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_1_MPORT_en & dataArray_27_1_MPORT_mask) begin
      dataArray_27_1[dataArray_27_1_MPORT_addr] <= dataArray_27_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_2_MPORT_en & dataArray_27_2_MPORT_mask) begin
      dataArray_27_2[dataArray_27_2_MPORT_addr] <= dataArray_27_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_3_MPORT_en & dataArray_27_3_MPORT_mask) begin
      dataArray_27_3[dataArray_27_3_MPORT_addr] <= dataArray_27_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_4_MPORT_en & dataArray_27_4_MPORT_mask) begin
      dataArray_27_4[dataArray_27_4_MPORT_addr] <= dataArray_27_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_5_MPORT_en & dataArray_27_5_MPORT_mask) begin
      dataArray_27_5[dataArray_27_5_MPORT_addr] <= dataArray_27_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_6_MPORT_en & dataArray_27_6_MPORT_mask) begin
      dataArray_27_6[dataArray_27_6_MPORT_addr] <= dataArray_27_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_7_MPORT_en & dataArray_27_7_MPORT_mask) begin
      dataArray_27_7[dataArray_27_7_MPORT_addr] <= dataArray_27_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_8_MPORT_en & dataArray_27_8_MPORT_mask) begin
      dataArray_27_8[dataArray_27_8_MPORT_addr] <= dataArray_27_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_9_MPORT_en & dataArray_27_9_MPORT_mask) begin
      dataArray_27_9[dataArray_27_9_MPORT_addr] <= dataArray_27_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_10_MPORT_en & dataArray_27_10_MPORT_mask) begin
      dataArray_27_10[dataArray_27_10_MPORT_addr] <= dataArray_27_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_11_MPORT_en & dataArray_27_11_MPORT_mask) begin
      dataArray_27_11[dataArray_27_11_MPORT_addr] <= dataArray_27_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_12_MPORT_en & dataArray_27_12_MPORT_mask) begin
      dataArray_27_12[dataArray_27_12_MPORT_addr] <= dataArray_27_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_13_MPORT_en & dataArray_27_13_MPORT_mask) begin
      dataArray_27_13[dataArray_27_13_MPORT_addr] <= dataArray_27_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_14_MPORT_en & dataArray_27_14_MPORT_mask) begin
      dataArray_27_14[dataArray_27_14_MPORT_addr] <= dataArray_27_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_27_15_MPORT_en & dataArray_27_15_MPORT_mask) begin
      dataArray_27_15[dataArray_27_15_MPORT_addr] <= dataArray_27_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_27_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_27_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_27_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_27_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_0_MPORT_en & dataArray_28_0_MPORT_mask) begin
      dataArray_28_0[dataArray_28_0_MPORT_addr] <= dataArray_28_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_1_MPORT_en & dataArray_28_1_MPORT_mask) begin
      dataArray_28_1[dataArray_28_1_MPORT_addr] <= dataArray_28_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_2_MPORT_en & dataArray_28_2_MPORT_mask) begin
      dataArray_28_2[dataArray_28_2_MPORT_addr] <= dataArray_28_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_3_MPORT_en & dataArray_28_3_MPORT_mask) begin
      dataArray_28_3[dataArray_28_3_MPORT_addr] <= dataArray_28_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_4_MPORT_en & dataArray_28_4_MPORT_mask) begin
      dataArray_28_4[dataArray_28_4_MPORT_addr] <= dataArray_28_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_5_MPORT_en & dataArray_28_5_MPORT_mask) begin
      dataArray_28_5[dataArray_28_5_MPORT_addr] <= dataArray_28_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_6_MPORT_en & dataArray_28_6_MPORT_mask) begin
      dataArray_28_6[dataArray_28_6_MPORT_addr] <= dataArray_28_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_7_MPORT_en & dataArray_28_7_MPORT_mask) begin
      dataArray_28_7[dataArray_28_7_MPORT_addr] <= dataArray_28_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_8_MPORT_en & dataArray_28_8_MPORT_mask) begin
      dataArray_28_8[dataArray_28_8_MPORT_addr] <= dataArray_28_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_9_MPORT_en & dataArray_28_9_MPORT_mask) begin
      dataArray_28_9[dataArray_28_9_MPORT_addr] <= dataArray_28_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_10_MPORT_en & dataArray_28_10_MPORT_mask) begin
      dataArray_28_10[dataArray_28_10_MPORT_addr] <= dataArray_28_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_11_MPORT_en & dataArray_28_11_MPORT_mask) begin
      dataArray_28_11[dataArray_28_11_MPORT_addr] <= dataArray_28_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_12_MPORT_en & dataArray_28_12_MPORT_mask) begin
      dataArray_28_12[dataArray_28_12_MPORT_addr] <= dataArray_28_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_13_MPORT_en & dataArray_28_13_MPORT_mask) begin
      dataArray_28_13[dataArray_28_13_MPORT_addr] <= dataArray_28_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_14_MPORT_en & dataArray_28_14_MPORT_mask) begin
      dataArray_28_14[dataArray_28_14_MPORT_addr] <= dataArray_28_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_28_15_MPORT_en & dataArray_28_15_MPORT_mask) begin
      dataArray_28_15[dataArray_28_15_MPORT_addr] <= dataArray_28_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_28_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_28_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_28_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_28_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_0_MPORT_en & dataArray_29_0_MPORT_mask) begin
      dataArray_29_0[dataArray_29_0_MPORT_addr] <= dataArray_29_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_1_MPORT_en & dataArray_29_1_MPORT_mask) begin
      dataArray_29_1[dataArray_29_1_MPORT_addr] <= dataArray_29_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_2_MPORT_en & dataArray_29_2_MPORT_mask) begin
      dataArray_29_2[dataArray_29_2_MPORT_addr] <= dataArray_29_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_3_MPORT_en & dataArray_29_3_MPORT_mask) begin
      dataArray_29_3[dataArray_29_3_MPORT_addr] <= dataArray_29_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_4_MPORT_en & dataArray_29_4_MPORT_mask) begin
      dataArray_29_4[dataArray_29_4_MPORT_addr] <= dataArray_29_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_5_MPORT_en & dataArray_29_5_MPORT_mask) begin
      dataArray_29_5[dataArray_29_5_MPORT_addr] <= dataArray_29_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_6_MPORT_en & dataArray_29_6_MPORT_mask) begin
      dataArray_29_6[dataArray_29_6_MPORT_addr] <= dataArray_29_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_7_MPORT_en & dataArray_29_7_MPORT_mask) begin
      dataArray_29_7[dataArray_29_7_MPORT_addr] <= dataArray_29_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_8_MPORT_en & dataArray_29_8_MPORT_mask) begin
      dataArray_29_8[dataArray_29_8_MPORT_addr] <= dataArray_29_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_9_MPORT_en & dataArray_29_9_MPORT_mask) begin
      dataArray_29_9[dataArray_29_9_MPORT_addr] <= dataArray_29_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_10_MPORT_en & dataArray_29_10_MPORT_mask) begin
      dataArray_29_10[dataArray_29_10_MPORT_addr] <= dataArray_29_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_11_MPORT_en & dataArray_29_11_MPORT_mask) begin
      dataArray_29_11[dataArray_29_11_MPORT_addr] <= dataArray_29_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_12_MPORT_en & dataArray_29_12_MPORT_mask) begin
      dataArray_29_12[dataArray_29_12_MPORT_addr] <= dataArray_29_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_13_MPORT_en & dataArray_29_13_MPORT_mask) begin
      dataArray_29_13[dataArray_29_13_MPORT_addr] <= dataArray_29_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_14_MPORT_en & dataArray_29_14_MPORT_mask) begin
      dataArray_29_14[dataArray_29_14_MPORT_addr] <= dataArray_29_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_29_15_MPORT_en & dataArray_29_15_MPORT_mask) begin
      dataArray_29_15[dataArray_29_15_MPORT_addr] <= dataArray_29_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_29_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_29_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_29_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_29_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_0_MPORT_en & dataArray_30_0_MPORT_mask) begin
      dataArray_30_0[dataArray_30_0_MPORT_addr] <= dataArray_30_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_1_MPORT_en & dataArray_30_1_MPORT_mask) begin
      dataArray_30_1[dataArray_30_1_MPORT_addr] <= dataArray_30_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_2_MPORT_en & dataArray_30_2_MPORT_mask) begin
      dataArray_30_2[dataArray_30_2_MPORT_addr] <= dataArray_30_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_3_MPORT_en & dataArray_30_3_MPORT_mask) begin
      dataArray_30_3[dataArray_30_3_MPORT_addr] <= dataArray_30_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_4_MPORT_en & dataArray_30_4_MPORT_mask) begin
      dataArray_30_4[dataArray_30_4_MPORT_addr] <= dataArray_30_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_5_MPORT_en & dataArray_30_5_MPORT_mask) begin
      dataArray_30_5[dataArray_30_5_MPORT_addr] <= dataArray_30_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_6_MPORT_en & dataArray_30_6_MPORT_mask) begin
      dataArray_30_6[dataArray_30_6_MPORT_addr] <= dataArray_30_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_7_MPORT_en & dataArray_30_7_MPORT_mask) begin
      dataArray_30_7[dataArray_30_7_MPORT_addr] <= dataArray_30_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_8_MPORT_en & dataArray_30_8_MPORT_mask) begin
      dataArray_30_8[dataArray_30_8_MPORT_addr] <= dataArray_30_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_9_MPORT_en & dataArray_30_9_MPORT_mask) begin
      dataArray_30_9[dataArray_30_9_MPORT_addr] <= dataArray_30_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_10_MPORT_en & dataArray_30_10_MPORT_mask) begin
      dataArray_30_10[dataArray_30_10_MPORT_addr] <= dataArray_30_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_11_MPORT_en & dataArray_30_11_MPORT_mask) begin
      dataArray_30_11[dataArray_30_11_MPORT_addr] <= dataArray_30_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_12_MPORT_en & dataArray_30_12_MPORT_mask) begin
      dataArray_30_12[dataArray_30_12_MPORT_addr] <= dataArray_30_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_13_MPORT_en & dataArray_30_13_MPORT_mask) begin
      dataArray_30_13[dataArray_30_13_MPORT_addr] <= dataArray_30_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_14_MPORT_en & dataArray_30_14_MPORT_mask) begin
      dataArray_30_14[dataArray_30_14_MPORT_addr] <= dataArray_30_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_30_15_MPORT_en & dataArray_30_15_MPORT_mask) begin
      dataArray_30_15[dataArray_30_15_MPORT_addr] <= dataArray_30_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_30_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_30_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_30_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_30_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_0_MPORT_en & dataArray_31_0_MPORT_mask) begin
      dataArray_31_0[dataArray_31_0_MPORT_addr] <= dataArray_31_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_1_MPORT_en & dataArray_31_1_MPORT_mask) begin
      dataArray_31_1[dataArray_31_1_MPORT_addr] <= dataArray_31_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_2_MPORT_en & dataArray_31_2_MPORT_mask) begin
      dataArray_31_2[dataArray_31_2_MPORT_addr] <= dataArray_31_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_3_MPORT_en & dataArray_31_3_MPORT_mask) begin
      dataArray_31_3[dataArray_31_3_MPORT_addr] <= dataArray_31_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_4_MPORT_en & dataArray_31_4_MPORT_mask) begin
      dataArray_31_4[dataArray_31_4_MPORT_addr] <= dataArray_31_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_5_MPORT_en & dataArray_31_5_MPORT_mask) begin
      dataArray_31_5[dataArray_31_5_MPORT_addr] <= dataArray_31_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_6_MPORT_en & dataArray_31_6_MPORT_mask) begin
      dataArray_31_6[dataArray_31_6_MPORT_addr] <= dataArray_31_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_7_MPORT_en & dataArray_31_7_MPORT_mask) begin
      dataArray_31_7[dataArray_31_7_MPORT_addr] <= dataArray_31_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_8_MPORT_en & dataArray_31_8_MPORT_mask) begin
      dataArray_31_8[dataArray_31_8_MPORT_addr] <= dataArray_31_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_9_MPORT_en & dataArray_31_9_MPORT_mask) begin
      dataArray_31_9[dataArray_31_9_MPORT_addr] <= dataArray_31_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_10_MPORT_en & dataArray_31_10_MPORT_mask) begin
      dataArray_31_10[dataArray_31_10_MPORT_addr] <= dataArray_31_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_11_MPORT_en & dataArray_31_11_MPORT_mask) begin
      dataArray_31_11[dataArray_31_11_MPORT_addr] <= dataArray_31_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_12_MPORT_en & dataArray_31_12_MPORT_mask) begin
      dataArray_31_12[dataArray_31_12_MPORT_addr] <= dataArray_31_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_13_MPORT_en & dataArray_31_13_MPORT_mask) begin
      dataArray_31_13[dataArray_31_13_MPORT_addr] <= dataArray_31_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_14_MPORT_en & dataArray_31_14_MPORT_mask) begin
      dataArray_31_14[dataArray_31_14_MPORT_addr] <= dataArray_31_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_31_15_MPORT_en & dataArray_31_15_MPORT_mask) begin
      dataArray_31_15[dataArray_31_15_MPORT_addr] <= dataArray_31_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_31_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_31_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_31_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_31_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_0_MPORT_en & dataArray_32_0_MPORT_mask) begin
      dataArray_32_0[dataArray_32_0_MPORT_addr] <= dataArray_32_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_1_MPORT_en & dataArray_32_1_MPORT_mask) begin
      dataArray_32_1[dataArray_32_1_MPORT_addr] <= dataArray_32_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_2_MPORT_en & dataArray_32_2_MPORT_mask) begin
      dataArray_32_2[dataArray_32_2_MPORT_addr] <= dataArray_32_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_3_MPORT_en & dataArray_32_3_MPORT_mask) begin
      dataArray_32_3[dataArray_32_3_MPORT_addr] <= dataArray_32_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_4_MPORT_en & dataArray_32_4_MPORT_mask) begin
      dataArray_32_4[dataArray_32_4_MPORT_addr] <= dataArray_32_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_5_MPORT_en & dataArray_32_5_MPORT_mask) begin
      dataArray_32_5[dataArray_32_5_MPORT_addr] <= dataArray_32_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_6_MPORT_en & dataArray_32_6_MPORT_mask) begin
      dataArray_32_6[dataArray_32_6_MPORT_addr] <= dataArray_32_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_7_MPORT_en & dataArray_32_7_MPORT_mask) begin
      dataArray_32_7[dataArray_32_7_MPORT_addr] <= dataArray_32_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_8_MPORT_en & dataArray_32_8_MPORT_mask) begin
      dataArray_32_8[dataArray_32_8_MPORT_addr] <= dataArray_32_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_9_MPORT_en & dataArray_32_9_MPORT_mask) begin
      dataArray_32_9[dataArray_32_9_MPORT_addr] <= dataArray_32_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_10_MPORT_en & dataArray_32_10_MPORT_mask) begin
      dataArray_32_10[dataArray_32_10_MPORT_addr] <= dataArray_32_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_11_MPORT_en & dataArray_32_11_MPORT_mask) begin
      dataArray_32_11[dataArray_32_11_MPORT_addr] <= dataArray_32_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_12_MPORT_en & dataArray_32_12_MPORT_mask) begin
      dataArray_32_12[dataArray_32_12_MPORT_addr] <= dataArray_32_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_13_MPORT_en & dataArray_32_13_MPORT_mask) begin
      dataArray_32_13[dataArray_32_13_MPORT_addr] <= dataArray_32_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_14_MPORT_en & dataArray_32_14_MPORT_mask) begin
      dataArray_32_14[dataArray_32_14_MPORT_addr] <= dataArray_32_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_32_15_MPORT_en & dataArray_32_15_MPORT_mask) begin
      dataArray_32_15[dataArray_32_15_MPORT_addr] <= dataArray_32_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_32_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_32_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_32_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_32_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_0_MPORT_en & dataArray_33_0_MPORT_mask) begin
      dataArray_33_0[dataArray_33_0_MPORT_addr] <= dataArray_33_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_1_MPORT_en & dataArray_33_1_MPORT_mask) begin
      dataArray_33_1[dataArray_33_1_MPORT_addr] <= dataArray_33_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_2_MPORT_en & dataArray_33_2_MPORT_mask) begin
      dataArray_33_2[dataArray_33_2_MPORT_addr] <= dataArray_33_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_3_MPORT_en & dataArray_33_3_MPORT_mask) begin
      dataArray_33_3[dataArray_33_3_MPORT_addr] <= dataArray_33_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_4_MPORT_en & dataArray_33_4_MPORT_mask) begin
      dataArray_33_4[dataArray_33_4_MPORT_addr] <= dataArray_33_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_5_MPORT_en & dataArray_33_5_MPORT_mask) begin
      dataArray_33_5[dataArray_33_5_MPORT_addr] <= dataArray_33_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_6_MPORT_en & dataArray_33_6_MPORT_mask) begin
      dataArray_33_6[dataArray_33_6_MPORT_addr] <= dataArray_33_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_7_MPORT_en & dataArray_33_7_MPORT_mask) begin
      dataArray_33_7[dataArray_33_7_MPORT_addr] <= dataArray_33_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_8_MPORT_en & dataArray_33_8_MPORT_mask) begin
      dataArray_33_8[dataArray_33_8_MPORT_addr] <= dataArray_33_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_9_MPORT_en & dataArray_33_9_MPORT_mask) begin
      dataArray_33_9[dataArray_33_9_MPORT_addr] <= dataArray_33_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_10_MPORT_en & dataArray_33_10_MPORT_mask) begin
      dataArray_33_10[dataArray_33_10_MPORT_addr] <= dataArray_33_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_11_MPORT_en & dataArray_33_11_MPORT_mask) begin
      dataArray_33_11[dataArray_33_11_MPORT_addr] <= dataArray_33_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_12_MPORT_en & dataArray_33_12_MPORT_mask) begin
      dataArray_33_12[dataArray_33_12_MPORT_addr] <= dataArray_33_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_13_MPORT_en & dataArray_33_13_MPORT_mask) begin
      dataArray_33_13[dataArray_33_13_MPORT_addr] <= dataArray_33_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_14_MPORT_en & dataArray_33_14_MPORT_mask) begin
      dataArray_33_14[dataArray_33_14_MPORT_addr] <= dataArray_33_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_33_15_MPORT_en & dataArray_33_15_MPORT_mask) begin
      dataArray_33_15[dataArray_33_15_MPORT_addr] <= dataArray_33_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_33_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_33_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_33_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_33_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_0_MPORT_en & dataArray_34_0_MPORT_mask) begin
      dataArray_34_0[dataArray_34_0_MPORT_addr] <= dataArray_34_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_1_MPORT_en & dataArray_34_1_MPORT_mask) begin
      dataArray_34_1[dataArray_34_1_MPORT_addr] <= dataArray_34_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_2_MPORT_en & dataArray_34_2_MPORT_mask) begin
      dataArray_34_2[dataArray_34_2_MPORT_addr] <= dataArray_34_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_3_MPORT_en & dataArray_34_3_MPORT_mask) begin
      dataArray_34_3[dataArray_34_3_MPORT_addr] <= dataArray_34_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_4_MPORT_en & dataArray_34_4_MPORT_mask) begin
      dataArray_34_4[dataArray_34_4_MPORT_addr] <= dataArray_34_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_5_MPORT_en & dataArray_34_5_MPORT_mask) begin
      dataArray_34_5[dataArray_34_5_MPORT_addr] <= dataArray_34_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_6_MPORT_en & dataArray_34_6_MPORT_mask) begin
      dataArray_34_6[dataArray_34_6_MPORT_addr] <= dataArray_34_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_7_MPORT_en & dataArray_34_7_MPORT_mask) begin
      dataArray_34_7[dataArray_34_7_MPORT_addr] <= dataArray_34_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_8_MPORT_en & dataArray_34_8_MPORT_mask) begin
      dataArray_34_8[dataArray_34_8_MPORT_addr] <= dataArray_34_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_9_MPORT_en & dataArray_34_9_MPORT_mask) begin
      dataArray_34_9[dataArray_34_9_MPORT_addr] <= dataArray_34_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_10_MPORT_en & dataArray_34_10_MPORT_mask) begin
      dataArray_34_10[dataArray_34_10_MPORT_addr] <= dataArray_34_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_11_MPORT_en & dataArray_34_11_MPORT_mask) begin
      dataArray_34_11[dataArray_34_11_MPORT_addr] <= dataArray_34_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_12_MPORT_en & dataArray_34_12_MPORT_mask) begin
      dataArray_34_12[dataArray_34_12_MPORT_addr] <= dataArray_34_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_13_MPORT_en & dataArray_34_13_MPORT_mask) begin
      dataArray_34_13[dataArray_34_13_MPORT_addr] <= dataArray_34_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_14_MPORT_en & dataArray_34_14_MPORT_mask) begin
      dataArray_34_14[dataArray_34_14_MPORT_addr] <= dataArray_34_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_34_15_MPORT_en & dataArray_34_15_MPORT_mask) begin
      dataArray_34_15[dataArray_34_15_MPORT_addr] <= dataArray_34_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_34_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_34_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_34_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_34_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_0_MPORT_en & dataArray_35_0_MPORT_mask) begin
      dataArray_35_0[dataArray_35_0_MPORT_addr] <= dataArray_35_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_1_MPORT_en & dataArray_35_1_MPORT_mask) begin
      dataArray_35_1[dataArray_35_1_MPORT_addr] <= dataArray_35_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_2_MPORT_en & dataArray_35_2_MPORT_mask) begin
      dataArray_35_2[dataArray_35_2_MPORT_addr] <= dataArray_35_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_3_MPORT_en & dataArray_35_3_MPORT_mask) begin
      dataArray_35_3[dataArray_35_3_MPORT_addr] <= dataArray_35_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_4_MPORT_en & dataArray_35_4_MPORT_mask) begin
      dataArray_35_4[dataArray_35_4_MPORT_addr] <= dataArray_35_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_5_MPORT_en & dataArray_35_5_MPORT_mask) begin
      dataArray_35_5[dataArray_35_5_MPORT_addr] <= dataArray_35_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_6_MPORT_en & dataArray_35_6_MPORT_mask) begin
      dataArray_35_6[dataArray_35_6_MPORT_addr] <= dataArray_35_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_7_MPORT_en & dataArray_35_7_MPORT_mask) begin
      dataArray_35_7[dataArray_35_7_MPORT_addr] <= dataArray_35_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_8_MPORT_en & dataArray_35_8_MPORT_mask) begin
      dataArray_35_8[dataArray_35_8_MPORT_addr] <= dataArray_35_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_9_MPORT_en & dataArray_35_9_MPORT_mask) begin
      dataArray_35_9[dataArray_35_9_MPORT_addr] <= dataArray_35_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_10_MPORT_en & dataArray_35_10_MPORT_mask) begin
      dataArray_35_10[dataArray_35_10_MPORT_addr] <= dataArray_35_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_11_MPORT_en & dataArray_35_11_MPORT_mask) begin
      dataArray_35_11[dataArray_35_11_MPORT_addr] <= dataArray_35_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_12_MPORT_en & dataArray_35_12_MPORT_mask) begin
      dataArray_35_12[dataArray_35_12_MPORT_addr] <= dataArray_35_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_13_MPORT_en & dataArray_35_13_MPORT_mask) begin
      dataArray_35_13[dataArray_35_13_MPORT_addr] <= dataArray_35_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_14_MPORT_en & dataArray_35_14_MPORT_mask) begin
      dataArray_35_14[dataArray_35_14_MPORT_addr] <= dataArray_35_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_35_15_MPORT_en & dataArray_35_15_MPORT_mask) begin
      dataArray_35_15[dataArray_35_15_MPORT_addr] <= dataArray_35_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_35_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_35_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_35_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_35_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_0_MPORT_en & dataArray_36_0_MPORT_mask) begin
      dataArray_36_0[dataArray_36_0_MPORT_addr] <= dataArray_36_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_1_MPORT_en & dataArray_36_1_MPORT_mask) begin
      dataArray_36_1[dataArray_36_1_MPORT_addr] <= dataArray_36_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_2_MPORT_en & dataArray_36_2_MPORT_mask) begin
      dataArray_36_2[dataArray_36_2_MPORT_addr] <= dataArray_36_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_3_MPORT_en & dataArray_36_3_MPORT_mask) begin
      dataArray_36_3[dataArray_36_3_MPORT_addr] <= dataArray_36_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_4_MPORT_en & dataArray_36_4_MPORT_mask) begin
      dataArray_36_4[dataArray_36_4_MPORT_addr] <= dataArray_36_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_5_MPORT_en & dataArray_36_5_MPORT_mask) begin
      dataArray_36_5[dataArray_36_5_MPORT_addr] <= dataArray_36_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_6_MPORT_en & dataArray_36_6_MPORT_mask) begin
      dataArray_36_6[dataArray_36_6_MPORT_addr] <= dataArray_36_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_7_MPORT_en & dataArray_36_7_MPORT_mask) begin
      dataArray_36_7[dataArray_36_7_MPORT_addr] <= dataArray_36_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_8_MPORT_en & dataArray_36_8_MPORT_mask) begin
      dataArray_36_8[dataArray_36_8_MPORT_addr] <= dataArray_36_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_9_MPORT_en & dataArray_36_9_MPORT_mask) begin
      dataArray_36_9[dataArray_36_9_MPORT_addr] <= dataArray_36_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_10_MPORT_en & dataArray_36_10_MPORT_mask) begin
      dataArray_36_10[dataArray_36_10_MPORT_addr] <= dataArray_36_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_11_MPORT_en & dataArray_36_11_MPORT_mask) begin
      dataArray_36_11[dataArray_36_11_MPORT_addr] <= dataArray_36_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_12_MPORT_en & dataArray_36_12_MPORT_mask) begin
      dataArray_36_12[dataArray_36_12_MPORT_addr] <= dataArray_36_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_13_MPORT_en & dataArray_36_13_MPORT_mask) begin
      dataArray_36_13[dataArray_36_13_MPORT_addr] <= dataArray_36_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_14_MPORT_en & dataArray_36_14_MPORT_mask) begin
      dataArray_36_14[dataArray_36_14_MPORT_addr] <= dataArray_36_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_36_15_MPORT_en & dataArray_36_15_MPORT_mask) begin
      dataArray_36_15[dataArray_36_15_MPORT_addr] <= dataArray_36_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_36_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_36_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_36_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_36_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_0_MPORT_en & dataArray_37_0_MPORT_mask) begin
      dataArray_37_0[dataArray_37_0_MPORT_addr] <= dataArray_37_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_1_MPORT_en & dataArray_37_1_MPORT_mask) begin
      dataArray_37_1[dataArray_37_1_MPORT_addr] <= dataArray_37_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_2_MPORT_en & dataArray_37_2_MPORT_mask) begin
      dataArray_37_2[dataArray_37_2_MPORT_addr] <= dataArray_37_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_3_MPORT_en & dataArray_37_3_MPORT_mask) begin
      dataArray_37_3[dataArray_37_3_MPORT_addr] <= dataArray_37_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_4_MPORT_en & dataArray_37_4_MPORT_mask) begin
      dataArray_37_4[dataArray_37_4_MPORT_addr] <= dataArray_37_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_5_MPORT_en & dataArray_37_5_MPORT_mask) begin
      dataArray_37_5[dataArray_37_5_MPORT_addr] <= dataArray_37_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_6_MPORT_en & dataArray_37_6_MPORT_mask) begin
      dataArray_37_6[dataArray_37_6_MPORT_addr] <= dataArray_37_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_7_MPORT_en & dataArray_37_7_MPORT_mask) begin
      dataArray_37_7[dataArray_37_7_MPORT_addr] <= dataArray_37_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_8_MPORT_en & dataArray_37_8_MPORT_mask) begin
      dataArray_37_8[dataArray_37_8_MPORT_addr] <= dataArray_37_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_9_MPORT_en & dataArray_37_9_MPORT_mask) begin
      dataArray_37_9[dataArray_37_9_MPORT_addr] <= dataArray_37_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_10_MPORT_en & dataArray_37_10_MPORT_mask) begin
      dataArray_37_10[dataArray_37_10_MPORT_addr] <= dataArray_37_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_11_MPORT_en & dataArray_37_11_MPORT_mask) begin
      dataArray_37_11[dataArray_37_11_MPORT_addr] <= dataArray_37_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_12_MPORT_en & dataArray_37_12_MPORT_mask) begin
      dataArray_37_12[dataArray_37_12_MPORT_addr] <= dataArray_37_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_13_MPORT_en & dataArray_37_13_MPORT_mask) begin
      dataArray_37_13[dataArray_37_13_MPORT_addr] <= dataArray_37_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_14_MPORT_en & dataArray_37_14_MPORT_mask) begin
      dataArray_37_14[dataArray_37_14_MPORT_addr] <= dataArray_37_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_37_15_MPORT_en & dataArray_37_15_MPORT_mask) begin
      dataArray_37_15[dataArray_37_15_MPORT_addr] <= dataArray_37_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_37_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_37_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_37_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_37_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_0_MPORT_en & dataArray_38_0_MPORT_mask) begin
      dataArray_38_0[dataArray_38_0_MPORT_addr] <= dataArray_38_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_1_MPORT_en & dataArray_38_1_MPORT_mask) begin
      dataArray_38_1[dataArray_38_1_MPORT_addr] <= dataArray_38_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_2_MPORT_en & dataArray_38_2_MPORT_mask) begin
      dataArray_38_2[dataArray_38_2_MPORT_addr] <= dataArray_38_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_3_MPORT_en & dataArray_38_3_MPORT_mask) begin
      dataArray_38_3[dataArray_38_3_MPORT_addr] <= dataArray_38_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_4_MPORT_en & dataArray_38_4_MPORT_mask) begin
      dataArray_38_4[dataArray_38_4_MPORT_addr] <= dataArray_38_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_5_MPORT_en & dataArray_38_5_MPORT_mask) begin
      dataArray_38_5[dataArray_38_5_MPORT_addr] <= dataArray_38_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_6_MPORT_en & dataArray_38_6_MPORT_mask) begin
      dataArray_38_6[dataArray_38_6_MPORT_addr] <= dataArray_38_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_7_MPORT_en & dataArray_38_7_MPORT_mask) begin
      dataArray_38_7[dataArray_38_7_MPORT_addr] <= dataArray_38_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_8_MPORT_en & dataArray_38_8_MPORT_mask) begin
      dataArray_38_8[dataArray_38_8_MPORT_addr] <= dataArray_38_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_9_MPORT_en & dataArray_38_9_MPORT_mask) begin
      dataArray_38_9[dataArray_38_9_MPORT_addr] <= dataArray_38_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_10_MPORT_en & dataArray_38_10_MPORT_mask) begin
      dataArray_38_10[dataArray_38_10_MPORT_addr] <= dataArray_38_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_11_MPORT_en & dataArray_38_11_MPORT_mask) begin
      dataArray_38_11[dataArray_38_11_MPORT_addr] <= dataArray_38_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_12_MPORT_en & dataArray_38_12_MPORT_mask) begin
      dataArray_38_12[dataArray_38_12_MPORT_addr] <= dataArray_38_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_13_MPORT_en & dataArray_38_13_MPORT_mask) begin
      dataArray_38_13[dataArray_38_13_MPORT_addr] <= dataArray_38_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_14_MPORT_en & dataArray_38_14_MPORT_mask) begin
      dataArray_38_14[dataArray_38_14_MPORT_addr] <= dataArray_38_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_38_15_MPORT_en & dataArray_38_15_MPORT_mask) begin
      dataArray_38_15[dataArray_38_15_MPORT_addr] <= dataArray_38_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_38_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_38_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_38_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_38_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_0_MPORT_en & dataArray_39_0_MPORT_mask) begin
      dataArray_39_0[dataArray_39_0_MPORT_addr] <= dataArray_39_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_1_MPORT_en & dataArray_39_1_MPORT_mask) begin
      dataArray_39_1[dataArray_39_1_MPORT_addr] <= dataArray_39_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_2_MPORT_en & dataArray_39_2_MPORT_mask) begin
      dataArray_39_2[dataArray_39_2_MPORT_addr] <= dataArray_39_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_3_MPORT_en & dataArray_39_3_MPORT_mask) begin
      dataArray_39_3[dataArray_39_3_MPORT_addr] <= dataArray_39_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_4_MPORT_en & dataArray_39_4_MPORT_mask) begin
      dataArray_39_4[dataArray_39_4_MPORT_addr] <= dataArray_39_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_5_MPORT_en & dataArray_39_5_MPORT_mask) begin
      dataArray_39_5[dataArray_39_5_MPORT_addr] <= dataArray_39_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_6_MPORT_en & dataArray_39_6_MPORT_mask) begin
      dataArray_39_6[dataArray_39_6_MPORT_addr] <= dataArray_39_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_7_MPORT_en & dataArray_39_7_MPORT_mask) begin
      dataArray_39_7[dataArray_39_7_MPORT_addr] <= dataArray_39_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_8_MPORT_en & dataArray_39_8_MPORT_mask) begin
      dataArray_39_8[dataArray_39_8_MPORT_addr] <= dataArray_39_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_9_MPORT_en & dataArray_39_9_MPORT_mask) begin
      dataArray_39_9[dataArray_39_9_MPORT_addr] <= dataArray_39_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_10_MPORT_en & dataArray_39_10_MPORT_mask) begin
      dataArray_39_10[dataArray_39_10_MPORT_addr] <= dataArray_39_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_11_MPORT_en & dataArray_39_11_MPORT_mask) begin
      dataArray_39_11[dataArray_39_11_MPORT_addr] <= dataArray_39_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_12_MPORT_en & dataArray_39_12_MPORT_mask) begin
      dataArray_39_12[dataArray_39_12_MPORT_addr] <= dataArray_39_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_13_MPORT_en & dataArray_39_13_MPORT_mask) begin
      dataArray_39_13[dataArray_39_13_MPORT_addr] <= dataArray_39_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_14_MPORT_en & dataArray_39_14_MPORT_mask) begin
      dataArray_39_14[dataArray_39_14_MPORT_addr] <= dataArray_39_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_39_15_MPORT_en & dataArray_39_15_MPORT_mask) begin
      dataArray_39_15[dataArray_39_15_MPORT_addr] <= dataArray_39_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_39_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_39_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_39_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_39_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_0_MPORT_en & dataArray_40_0_MPORT_mask) begin
      dataArray_40_0[dataArray_40_0_MPORT_addr] <= dataArray_40_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_1_MPORT_en & dataArray_40_1_MPORT_mask) begin
      dataArray_40_1[dataArray_40_1_MPORT_addr] <= dataArray_40_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_2_MPORT_en & dataArray_40_2_MPORT_mask) begin
      dataArray_40_2[dataArray_40_2_MPORT_addr] <= dataArray_40_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_3_MPORT_en & dataArray_40_3_MPORT_mask) begin
      dataArray_40_3[dataArray_40_3_MPORT_addr] <= dataArray_40_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_4_MPORT_en & dataArray_40_4_MPORT_mask) begin
      dataArray_40_4[dataArray_40_4_MPORT_addr] <= dataArray_40_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_5_MPORT_en & dataArray_40_5_MPORT_mask) begin
      dataArray_40_5[dataArray_40_5_MPORT_addr] <= dataArray_40_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_6_MPORT_en & dataArray_40_6_MPORT_mask) begin
      dataArray_40_6[dataArray_40_6_MPORT_addr] <= dataArray_40_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_7_MPORT_en & dataArray_40_7_MPORT_mask) begin
      dataArray_40_7[dataArray_40_7_MPORT_addr] <= dataArray_40_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_8_MPORT_en & dataArray_40_8_MPORT_mask) begin
      dataArray_40_8[dataArray_40_8_MPORT_addr] <= dataArray_40_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_9_MPORT_en & dataArray_40_9_MPORT_mask) begin
      dataArray_40_9[dataArray_40_9_MPORT_addr] <= dataArray_40_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_10_MPORT_en & dataArray_40_10_MPORT_mask) begin
      dataArray_40_10[dataArray_40_10_MPORT_addr] <= dataArray_40_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_11_MPORT_en & dataArray_40_11_MPORT_mask) begin
      dataArray_40_11[dataArray_40_11_MPORT_addr] <= dataArray_40_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_12_MPORT_en & dataArray_40_12_MPORT_mask) begin
      dataArray_40_12[dataArray_40_12_MPORT_addr] <= dataArray_40_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_13_MPORT_en & dataArray_40_13_MPORT_mask) begin
      dataArray_40_13[dataArray_40_13_MPORT_addr] <= dataArray_40_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_14_MPORT_en & dataArray_40_14_MPORT_mask) begin
      dataArray_40_14[dataArray_40_14_MPORT_addr] <= dataArray_40_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_40_15_MPORT_en & dataArray_40_15_MPORT_mask) begin
      dataArray_40_15[dataArray_40_15_MPORT_addr] <= dataArray_40_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_40_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_40_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_40_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_40_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_0_MPORT_en & dataArray_41_0_MPORT_mask) begin
      dataArray_41_0[dataArray_41_0_MPORT_addr] <= dataArray_41_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_1_MPORT_en & dataArray_41_1_MPORT_mask) begin
      dataArray_41_1[dataArray_41_1_MPORT_addr] <= dataArray_41_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_2_MPORT_en & dataArray_41_2_MPORT_mask) begin
      dataArray_41_2[dataArray_41_2_MPORT_addr] <= dataArray_41_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_3_MPORT_en & dataArray_41_3_MPORT_mask) begin
      dataArray_41_3[dataArray_41_3_MPORT_addr] <= dataArray_41_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_4_MPORT_en & dataArray_41_4_MPORT_mask) begin
      dataArray_41_4[dataArray_41_4_MPORT_addr] <= dataArray_41_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_5_MPORT_en & dataArray_41_5_MPORT_mask) begin
      dataArray_41_5[dataArray_41_5_MPORT_addr] <= dataArray_41_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_6_MPORT_en & dataArray_41_6_MPORT_mask) begin
      dataArray_41_6[dataArray_41_6_MPORT_addr] <= dataArray_41_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_7_MPORT_en & dataArray_41_7_MPORT_mask) begin
      dataArray_41_7[dataArray_41_7_MPORT_addr] <= dataArray_41_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_8_MPORT_en & dataArray_41_8_MPORT_mask) begin
      dataArray_41_8[dataArray_41_8_MPORT_addr] <= dataArray_41_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_9_MPORT_en & dataArray_41_9_MPORT_mask) begin
      dataArray_41_9[dataArray_41_9_MPORT_addr] <= dataArray_41_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_10_MPORT_en & dataArray_41_10_MPORT_mask) begin
      dataArray_41_10[dataArray_41_10_MPORT_addr] <= dataArray_41_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_11_MPORT_en & dataArray_41_11_MPORT_mask) begin
      dataArray_41_11[dataArray_41_11_MPORT_addr] <= dataArray_41_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_12_MPORT_en & dataArray_41_12_MPORT_mask) begin
      dataArray_41_12[dataArray_41_12_MPORT_addr] <= dataArray_41_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_13_MPORT_en & dataArray_41_13_MPORT_mask) begin
      dataArray_41_13[dataArray_41_13_MPORT_addr] <= dataArray_41_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_14_MPORT_en & dataArray_41_14_MPORT_mask) begin
      dataArray_41_14[dataArray_41_14_MPORT_addr] <= dataArray_41_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_41_15_MPORT_en & dataArray_41_15_MPORT_mask) begin
      dataArray_41_15[dataArray_41_15_MPORT_addr] <= dataArray_41_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_41_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_41_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_41_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_41_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_0_MPORT_en & dataArray_42_0_MPORT_mask) begin
      dataArray_42_0[dataArray_42_0_MPORT_addr] <= dataArray_42_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_1_MPORT_en & dataArray_42_1_MPORT_mask) begin
      dataArray_42_1[dataArray_42_1_MPORT_addr] <= dataArray_42_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_2_MPORT_en & dataArray_42_2_MPORT_mask) begin
      dataArray_42_2[dataArray_42_2_MPORT_addr] <= dataArray_42_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_3_MPORT_en & dataArray_42_3_MPORT_mask) begin
      dataArray_42_3[dataArray_42_3_MPORT_addr] <= dataArray_42_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_4_MPORT_en & dataArray_42_4_MPORT_mask) begin
      dataArray_42_4[dataArray_42_4_MPORT_addr] <= dataArray_42_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_5_MPORT_en & dataArray_42_5_MPORT_mask) begin
      dataArray_42_5[dataArray_42_5_MPORT_addr] <= dataArray_42_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_6_MPORT_en & dataArray_42_6_MPORT_mask) begin
      dataArray_42_6[dataArray_42_6_MPORT_addr] <= dataArray_42_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_7_MPORT_en & dataArray_42_7_MPORT_mask) begin
      dataArray_42_7[dataArray_42_7_MPORT_addr] <= dataArray_42_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_8_MPORT_en & dataArray_42_8_MPORT_mask) begin
      dataArray_42_8[dataArray_42_8_MPORT_addr] <= dataArray_42_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_9_MPORT_en & dataArray_42_9_MPORT_mask) begin
      dataArray_42_9[dataArray_42_9_MPORT_addr] <= dataArray_42_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_10_MPORT_en & dataArray_42_10_MPORT_mask) begin
      dataArray_42_10[dataArray_42_10_MPORT_addr] <= dataArray_42_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_11_MPORT_en & dataArray_42_11_MPORT_mask) begin
      dataArray_42_11[dataArray_42_11_MPORT_addr] <= dataArray_42_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_12_MPORT_en & dataArray_42_12_MPORT_mask) begin
      dataArray_42_12[dataArray_42_12_MPORT_addr] <= dataArray_42_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_13_MPORT_en & dataArray_42_13_MPORT_mask) begin
      dataArray_42_13[dataArray_42_13_MPORT_addr] <= dataArray_42_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_14_MPORT_en & dataArray_42_14_MPORT_mask) begin
      dataArray_42_14[dataArray_42_14_MPORT_addr] <= dataArray_42_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_42_15_MPORT_en & dataArray_42_15_MPORT_mask) begin
      dataArray_42_15[dataArray_42_15_MPORT_addr] <= dataArray_42_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_42_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_42_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_42_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_42_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_0_MPORT_en & dataArray_43_0_MPORT_mask) begin
      dataArray_43_0[dataArray_43_0_MPORT_addr] <= dataArray_43_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_1_MPORT_en & dataArray_43_1_MPORT_mask) begin
      dataArray_43_1[dataArray_43_1_MPORT_addr] <= dataArray_43_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_2_MPORT_en & dataArray_43_2_MPORT_mask) begin
      dataArray_43_2[dataArray_43_2_MPORT_addr] <= dataArray_43_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_3_MPORT_en & dataArray_43_3_MPORT_mask) begin
      dataArray_43_3[dataArray_43_3_MPORT_addr] <= dataArray_43_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_4_MPORT_en & dataArray_43_4_MPORT_mask) begin
      dataArray_43_4[dataArray_43_4_MPORT_addr] <= dataArray_43_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_5_MPORT_en & dataArray_43_5_MPORT_mask) begin
      dataArray_43_5[dataArray_43_5_MPORT_addr] <= dataArray_43_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_6_MPORT_en & dataArray_43_6_MPORT_mask) begin
      dataArray_43_6[dataArray_43_6_MPORT_addr] <= dataArray_43_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_7_MPORT_en & dataArray_43_7_MPORT_mask) begin
      dataArray_43_7[dataArray_43_7_MPORT_addr] <= dataArray_43_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_8_MPORT_en & dataArray_43_8_MPORT_mask) begin
      dataArray_43_8[dataArray_43_8_MPORT_addr] <= dataArray_43_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_9_MPORT_en & dataArray_43_9_MPORT_mask) begin
      dataArray_43_9[dataArray_43_9_MPORT_addr] <= dataArray_43_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_10_MPORT_en & dataArray_43_10_MPORT_mask) begin
      dataArray_43_10[dataArray_43_10_MPORT_addr] <= dataArray_43_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_11_MPORT_en & dataArray_43_11_MPORT_mask) begin
      dataArray_43_11[dataArray_43_11_MPORT_addr] <= dataArray_43_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_12_MPORT_en & dataArray_43_12_MPORT_mask) begin
      dataArray_43_12[dataArray_43_12_MPORT_addr] <= dataArray_43_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_13_MPORT_en & dataArray_43_13_MPORT_mask) begin
      dataArray_43_13[dataArray_43_13_MPORT_addr] <= dataArray_43_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_14_MPORT_en & dataArray_43_14_MPORT_mask) begin
      dataArray_43_14[dataArray_43_14_MPORT_addr] <= dataArray_43_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_43_15_MPORT_en & dataArray_43_15_MPORT_mask) begin
      dataArray_43_15[dataArray_43_15_MPORT_addr] <= dataArray_43_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_43_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_43_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_43_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_43_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_0_MPORT_en & dataArray_44_0_MPORT_mask) begin
      dataArray_44_0[dataArray_44_0_MPORT_addr] <= dataArray_44_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_1_MPORT_en & dataArray_44_1_MPORT_mask) begin
      dataArray_44_1[dataArray_44_1_MPORT_addr] <= dataArray_44_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_2_MPORT_en & dataArray_44_2_MPORT_mask) begin
      dataArray_44_2[dataArray_44_2_MPORT_addr] <= dataArray_44_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_3_MPORT_en & dataArray_44_3_MPORT_mask) begin
      dataArray_44_3[dataArray_44_3_MPORT_addr] <= dataArray_44_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_4_MPORT_en & dataArray_44_4_MPORT_mask) begin
      dataArray_44_4[dataArray_44_4_MPORT_addr] <= dataArray_44_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_5_MPORT_en & dataArray_44_5_MPORT_mask) begin
      dataArray_44_5[dataArray_44_5_MPORT_addr] <= dataArray_44_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_6_MPORT_en & dataArray_44_6_MPORT_mask) begin
      dataArray_44_6[dataArray_44_6_MPORT_addr] <= dataArray_44_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_7_MPORT_en & dataArray_44_7_MPORT_mask) begin
      dataArray_44_7[dataArray_44_7_MPORT_addr] <= dataArray_44_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_8_MPORT_en & dataArray_44_8_MPORT_mask) begin
      dataArray_44_8[dataArray_44_8_MPORT_addr] <= dataArray_44_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_9_MPORT_en & dataArray_44_9_MPORT_mask) begin
      dataArray_44_9[dataArray_44_9_MPORT_addr] <= dataArray_44_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_10_MPORT_en & dataArray_44_10_MPORT_mask) begin
      dataArray_44_10[dataArray_44_10_MPORT_addr] <= dataArray_44_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_11_MPORT_en & dataArray_44_11_MPORT_mask) begin
      dataArray_44_11[dataArray_44_11_MPORT_addr] <= dataArray_44_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_12_MPORT_en & dataArray_44_12_MPORT_mask) begin
      dataArray_44_12[dataArray_44_12_MPORT_addr] <= dataArray_44_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_13_MPORT_en & dataArray_44_13_MPORT_mask) begin
      dataArray_44_13[dataArray_44_13_MPORT_addr] <= dataArray_44_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_14_MPORT_en & dataArray_44_14_MPORT_mask) begin
      dataArray_44_14[dataArray_44_14_MPORT_addr] <= dataArray_44_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_44_15_MPORT_en & dataArray_44_15_MPORT_mask) begin
      dataArray_44_15[dataArray_44_15_MPORT_addr] <= dataArray_44_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_44_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_44_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_44_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_44_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_0_MPORT_en & dataArray_45_0_MPORT_mask) begin
      dataArray_45_0[dataArray_45_0_MPORT_addr] <= dataArray_45_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_1_MPORT_en & dataArray_45_1_MPORT_mask) begin
      dataArray_45_1[dataArray_45_1_MPORT_addr] <= dataArray_45_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_2_MPORT_en & dataArray_45_2_MPORT_mask) begin
      dataArray_45_2[dataArray_45_2_MPORT_addr] <= dataArray_45_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_3_MPORT_en & dataArray_45_3_MPORT_mask) begin
      dataArray_45_3[dataArray_45_3_MPORT_addr] <= dataArray_45_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_4_MPORT_en & dataArray_45_4_MPORT_mask) begin
      dataArray_45_4[dataArray_45_4_MPORT_addr] <= dataArray_45_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_5_MPORT_en & dataArray_45_5_MPORT_mask) begin
      dataArray_45_5[dataArray_45_5_MPORT_addr] <= dataArray_45_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_6_MPORT_en & dataArray_45_6_MPORT_mask) begin
      dataArray_45_6[dataArray_45_6_MPORT_addr] <= dataArray_45_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_7_MPORT_en & dataArray_45_7_MPORT_mask) begin
      dataArray_45_7[dataArray_45_7_MPORT_addr] <= dataArray_45_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_8_MPORT_en & dataArray_45_8_MPORT_mask) begin
      dataArray_45_8[dataArray_45_8_MPORT_addr] <= dataArray_45_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_9_MPORT_en & dataArray_45_9_MPORT_mask) begin
      dataArray_45_9[dataArray_45_9_MPORT_addr] <= dataArray_45_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_10_MPORT_en & dataArray_45_10_MPORT_mask) begin
      dataArray_45_10[dataArray_45_10_MPORT_addr] <= dataArray_45_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_11_MPORT_en & dataArray_45_11_MPORT_mask) begin
      dataArray_45_11[dataArray_45_11_MPORT_addr] <= dataArray_45_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_12_MPORT_en & dataArray_45_12_MPORT_mask) begin
      dataArray_45_12[dataArray_45_12_MPORT_addr] <= dataArray_45_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_13_MPORT_en & dataArray_45_13_MPORT_mask) begin
      dataArray_45_13[dataArray_45_13_MPORT_addr] <= dataArray_45_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_14_MPORT_en & dataArray_45_14_MPORT_mask) begin
      dataArray_45_14[dataArray_45_14_MPORT_addr] <= dataArray_45_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_45_15_MPORT_en & dataArray_45_15_MPORT_mask) begin
      dataArray_45_15[dataArray_45_15_MPORT_addr] <= dataArray_45_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_45_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_45_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_45_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_45_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_0_MPORT_en & dataArray_46_0_MPORT_mask) begin
      dataArray_46_0[dataArray_46_0_MPORT_addr] <= dataArray_46_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_1_MPORT_en & dataArray_46_1_MPORT_mask) begin
      dataArray_46_1[dataArray_46_1_MPORT_addr] <= dataArray_46_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_2_MPORT_en & dataArray_46_2_MPORT_mask) begin
      dataArray_46_2[dataArray_46_2_MPORT_addr] <= dataArray_46_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_3_MPORT_en & dataArray_46_3_MPORT_mask) begin
      dataArray_46_3[dataArray_46_3_MPORT_addr] <= dataArray_46_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_4_MPORT_en & dataArray_46_4_MPORT_mask) begin
      dataArray_46_4[dataArray_46_4_MPORT_addr] <= dataArray_46_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_5_MPORT_en & dataArray_46_5_MPORT_mask) begin
      dataArray_46_5[dataArray_46_5_MPORT_addr] <= dataArray_46_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_6_MPORT_en & dataArray_46_6_MPORT_mask) begin
      dataArray_46_6[dataArray_46_6_MPORT_addr] <= dataArray_46_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_7_MPORT_en & dataArray_46_7_MPORT_mask) begin
      dataArray_46_7[dataArray_46_7_MPORT_addr] <= dataArray_46_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_8_MPORT_en & dataArray_46_8_MPORT_mask) begin
      dataArray_46_8[dataArray_46_8_MPORT_addr] <= dataArray_46_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_9_MPORT_en & dataArray_46_9_MPORT_mask) begin
      dataArray_46_9[dataArray_46_9_MPORT_addr] <= dataArray_46_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_10_MPORT_en & dataArray_46_10_MPORT_mask) begin
      dataArray_46_10[dataArray_46_10_MPORT_addr] <= dataArray_46_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_11_MPORT_en & dataArray_46_11_MPORT_mask) begin
      dataArray_46_11[dataArray_46_11_MPORT_addr] <= dataArray_46_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_12_MPORT_en & dataArray_46_12_MPORT_mask) begin
      dataArray_46_12[dataArray_46_12_MPORT_addr] <= dataArray_46_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_13_MPORT_en & dataArray_46_13_MPORT_mask) begin
      dataArray_46_13[dataArray_46_13_MPORT_addr] <= dataArray_46_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_14_MPORT_en & dataArray_46_14_MPORT_mask) begin
      dataArray_46_14[dataArray_46_14_MPORT_addr] <= dataArray_46_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_46_15_MPORT_en & dataArray_46_15_MPORT_mask) begin
      dataArray_46_15[dataArray_46_15_MPORT_addr] <= dataArray_46_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_46_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_46_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_46_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_46_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_0_MPORT_en & dataArray_47_0_MPORT_mask) begin
      dataArray_47_0[dataArray_47_0_MPORT_addr] <= dataArray_47_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_1_MPORT_en & dataArray_47_1_MPORT_mask) begin
      dataArray_47_1[dataArray_47_1_MPORT_addr] <= dataArray_47_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_2_MPORT_en & dataArray_47_2_MPORT_mask) begin
      dataArray_47_2[dataArray_47_2_MPORT_addr] <= dataArray_47_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_3_MPORT_en & dataArray_47_3_MPORT_mask) begin
      dataArray_47_3[dataArray_47_3_MPORT_addr] <= dataArray_47_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_4_MPORT_en & dataArray_47_4_MPORT_mask) begin
      dataArray_47_4[dataArray_47_4_MPORT_addr] <= dataArray_47_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_5_MPORT_en & dataArray_47_5_MPORT_mask) begin
      dataArray_47_5[dataArray_47_5_MPORT_addr] <= dataArray_47_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_6_MPORT_en & dataArray_47_6_MPORT_mask) begin
      dataArray_47_6[dataArray_47_6_MPORT_addr] <= dataArray_47_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_7_MPORT_en & dataArray_47_7_MPORT_mask) begin
      dataArray_47_7[dataArray_47_7_MPORT_addr] <= dataArray_47_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_8_MPORT_en & dataArray_47_8_MPORT_mask) begin
      dataArray_47_8[dataArray_47_8_MPORT_addr] <= dataArray_47_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_9_MPORT_en & dataArray_47_9_MPORT_mask) begin
      dataArray_47_9[dataArray_47_9_MPORT_addr] <= dataArray_47_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_10_MPORT_en & dataArray_47_10_MPORT_mask) begin
      dataArray_47_10[dataArray_47_10_MPORT_addr] <= dataArray_47_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_11_MPORT_en & dataArray_47_11_MPORT_mask) begin
      dataArray_47_11[dataArray_47_11_MPORT_addr] <= dataArray_47_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_12_MPORT_en & dataArray_47_12_MPORT_mask) begin
      dataArray_47_12[dataArray_47_12_MPORT_addr] <= dataArray_47_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_13_MPORT_en & dataArray_47_13_MPORT_mask) begin
      dataArray_47_13[dataArray_47_13_MPORT_addr] <= dataArray_47_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_14_MPORT_en & dataArray_47_14_MPORT_mask) begin
      dataArray_47_14[dataArray_47_14_MPORT_addr] <= dataArray_47_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_47_15_MPORT_en & dataArray_47_15_MPORT_mask) begin
      dataArray_47_15[dataArray_47_15_MPORT_addr] <= dataArray_47_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_47_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_47_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_47_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_47_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_0_MPORT_en & dataArray_48_0_MPORT_mask) begin
      dataArray_48_0[dataArray_48_0_MPORT_addr] <= dataArray_48_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_1_MPORT_en & dataArray_48_1_MPORT_mask) begin
      dataArray_48_1[dataArray_48_1_MPORT_addr] <= dataArray_48_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_2_MPORT_en & dataArray_48_2_MPORT_mask) begin
      dataArray_48_2[dataArray_48_2_MPORT_addr] <= dataArray_48_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_3_MPORT_en & dataArray_48_3_MPORT_mask) begin
      dataArray_48_3[dataArray_48_3_MPORT_addr] <= dataArray_48_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_4_MPORT_en & dataArray_48_4_MPORT_mask) begin
      dataArray_48_4[dataArray_48_4_MPORT_addr] <= dataArray_48_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_5_MPORT_en & dataArray_48_5_MPORT_mask) begin
      dataArray_48_5[dataArray_48_5_MPORT_addr] <= dataArray_48_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_6_MPORT_en & dataArray_48_6_MPORT_mask) begin
      dataArray_48_6[dataArray_48_6_MPORT_addr] <= dataArray_48_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_7_MPORT_en & dataArray_48_7_MPORT_mask) begin
      dataArray_48_7[dataArray_48_7_MPORT_addr] <= dataArray_48_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_8_MPORT_en & dataArray_48_8_MPORT_mask) begin
      dataArray_48_8[dataArray_48_8_MPORT_addr] <= dataArray_48_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_9_MPORT_en & dataArray_48_9_MPORT_mask) begin
      dataArray_48_9[dataArray_48_9_MPORT_addr] <= dataArray_48_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_10_MPORT_en & dataArray_48_10_MPORT_mask) begin
      dataArray_48_10[dataArray_48_10_MPORT_addr] <= dataArray_48_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_11_MPORT_en & dataArray_48_11_MPORT_mask) begin
      dataArray_48_11[dataArray_48_11_MPORT_addr] <= dataArray_48_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_12_MPORT_en & dataArray_48_12_MPORT_mask) begin
      dataArray_48_12[dataArray_48_12_MPORT_addr] <= dataArray_48_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_13_MPORT_en & dataArray_48_13_MPORT_mask) begin
      dataArray_48_13[dataArray_48_13_MPORT_addr] <= dataArray_48_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_14_MPORT_en & dataArray_48_14_MPORT_mask) begin
      dataArray_48_14[dataArray_48_14_MPORT_addr] <= dataArray_48_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_48_15_MPORT_en & dataArray_48_15_MPORT_mask) begin
      dataArray_48_15[dataArray_48_15_MPORT_addr] <= dataArray_48_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_48_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_48_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_48_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_48_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_0_MPORT_en & dataArray_49_0_MPORT_mask) begin
      dataArray_49_0[dataArray_49_0_MPORT_addr] <= dataArray_49_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_1_MPORT_en & dataArray_49_1_MPORT_mask) begin
      dataArray_49_1[dataArray_49_1_MPORT_addr] <= dataArray_49_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_2_MPORT_en & dataArray_49_2_MPORT_mask) begin
      dataArray_49_2[dataArray_49_2_MPORT_addr] <= dataArray_49_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_3_MPORT_en & dataArray_49_3_MPORT_mask) begin
      dataArray_49_3[dataArray_49_3_MPORT_addr] <= dataArray_49_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_4_MPORT_en & dataArray_49_4_MPORT_mask) begin
      dataArray_49_4[dataArray_49_4_MPORT_addr] <= dataArray_49_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_5_MPORT_en & dataArray_49_5_MPORT_mask) begin
      dataArray_49_5[dataArray_49_5_MPORT_addr] <= dataArray_49_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_6_MPORT_en & dataArray_49_6_MPORT_mask) begin
      dataArray_49_6[dataArray_49_6_MPORT_addr] <= dataArray_49_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_7_MPORT_en & dataArray_49_7_MPORT_mask) begin
      dataArray_49_7[dataArray_49_7_MPORT_addr] <= dataArray_49_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_8_MPORT_en & dataArray_49_8_MPORT_mask) begin
      dataArray_49_8[dataArray_49_8_MPORT_addr] <= dataArray_49_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_9_MPORT_en & dataArray_49_9_MPORT_mask) begin
      dataArray_49_9[dataArray_49_9_MPORT_addr] <= dataArray_49_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_10_MPORT_en & dataArray_49_10_MPORT_mask) begin
      dataArray_49_10[dataArray_49_10_MPORT_addr] <= dataArray_49_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_11_MPORT_en & dataArray_49_11_MPORT_mask) begin
      dataArray_49_11[dataArray_49_11_MPORT_addr] <= dataArray_49_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_12_MPORT_en & dataArray_49_12_MPORT_mask) begin
      dataArray_49_12[dataArray_49_12_MPORT_addr] <= dataArray_49_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_13_MPORT_en & dataArray_49_13_MPORT_mask) begin
      dataArray_49_13[dataArray_49_13_MPORT_addr] <= dataArray_49_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_14_MPORT_en & dataArray_49_14_MPORT_mask) begin
      dataArray_49_14[dataArray_49_14_MPORT_addr] <= dataArray_49_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_49_15_MPORT_en & dataArray_49_15_MPORT_mask) begin
      dataArray_49_15[dataArray_49_15_MPORT_addr] <= dataArray_49_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_49_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_49_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_49_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_49_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_0_MPORT_en & dataArray_50_0_MPORT_mask) begin
      dataArray_50_0[dataArray_50_0_MPORT_addr] <= dataArray_50_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_1_MPORT_en & dataArray_50_1_MPORT_mask) begin
      dataArray_50_1[dataArray_50_1_MPORT_addr] <= dataArray_50_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_2_MPORT_en & dataArray_50_2_MPORT_mask) begin
      dataArray_50_2[dataArray_50_2_MPORT_addr] <= dataArray_50_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_3_MPORT_en & dataArray_50_3_MPORT_mask) begin
      dataArray_50_3[dataArray_50_3_MPORT_addr] <= dataArray_50_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_4_MPORT_en & dataArray_50_4_MPORT_mask) begin
      dataArray_50_4[dataArray_50_4_MPORT_addr] <= dataArray_50_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_5_MPORT_en & dataArray_50_5_MPORT_mask) begin
      dataArray_50_5[dataArray_50_5_MPORT_addr] <= dataArray_50_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_6_MPORT_en & dataArray_50_6_MPORT_mask) begin
      dataArray_50_6[dataArray_50_6_MPORT_addr] <= dataArray_50_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_7_MPORT_en & dataArray_50_7_MPORT_mask) begin
      dataArray_50_7[dataArray_50_7_MPORT_addr] <= dataArray_50_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_8_MPORT_en & dataArray_50_8_MPORT_mask) begin
      dataArray_50_8[dataArray_50_8_MPORT_addr] <= dataArray_50_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_9_MPORT_en & dataArray_50_9_MPORT_mask) begin
      dataArray_50_9[dataArray_50_9_MPORT_addr] <= dataArray_50_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_10_MPORT_en & dataArray_50_10_MPORT_mask) begin
      dataArray_50_10[dataArray_50_10_MPORT_addr] <= dataArray_50_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_11_MPORT_en & dataArray_50_11_MPORT_mask) begin
      dataArray_50_11[dataArray_50_11_MPORT_addr] <= dataArray_50_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_12_MPORT_en & dataArray_50_12_MPORT_mask) begin
      dataArray_50_12[dataArray_50_12_MPORT_addr] <= dataArray_50_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_13_MPORT_en & dataArray_50_13_MPORT_mask) begin
      dataArray_50_13[dataArray_50_13_MPORT_addr] <= dataArray_50_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_14_MPORT_en & dataArray_50_14_MPORT_mask) begin
      dataArray_50_14[dataArray_50_14_MPORT_addr] <= dataArray_50_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_50_15_MPORT_en & dataArray_50_15_MPORT_mask) begin
      dataArray_50_15[dataArray_50_15_MPORT_addr] <= dataArray_50_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_50_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_50_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_50_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_50_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_0_MPORT_en & dataArray_51_0_MPORT_mask) begin
      dataArray_51_0[dataArray_51_0_MPORT_addr] <= dataArray_51_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_1_MPORT_en & dataArray_51_1_MPORT_mask) begin
      dataArray_51_1[dataArray_51_1_MPORT_addr] <= dataArray_51_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_2_MPORT_en & dataArray_51_2_MPORT_mask) begin
      dataArray_51_2[dataArray_51_2_MPORT_addr] <= dataArray_51_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_3_MPORT_en & dataArray_51_3_MPORT_mask) begin
      dataArray_51_3[dataArray_51_3_MPORT_addr] <= dataArray_51_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_4_MPORT_en & dataArray_51_4_MPORT_mask) begin
      dataArray_51_4[dataArray_51_4_MPORT_addr] <= dataArray_51_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_5_MPORT_en & dataArray_51_5_MPORT_mask) begin
      dataArray_51_5[dataArray_51_5_MPORT_addr] <= dataArray_51_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_6_MPORT_en & dataArray_51_6_MPORT_mask) begin
      dataArray_51_6[dataArray_51_6_MPORT_addr] <= dataArray_51_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_7_MPORT_en & dataArray_51_7_MPORT_mask) begin
      dataArray_51_7[dataArray_51_7_MPORT_addr] <= dataArray_51_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_8_MPORT_en & dataArray_51_8_MPORT_mask) begin
      dataArray_51_8[dataArray_51_8_MPORT_addr] <= dataArray_51_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_9_MPORT_en & dataArray_51_9_MPORT_mask) begin
      dataArray_51_9[dataArray_51_9_MPORT_addr] <= dataArray_51_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_10_MPORT_en & dataArray_51_10_MPORT_mask) begin
      dataArray_51_10[dataArray_51_10_MPORT_addr] <= dataArray_51_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_11_MPORT_en & dataArray_51_11_MPORT_mask) begin
      dataArray_51_11[dataArray_51_11_MPORT_addr] <= dataArray_51_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_12_MPORT_en & dataArray_51_12_MPORT_mask) begin
      dataArray_51_12[dataArray_51_12_MPORT_addr] <= dataArray_51_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_13_MPORT_en & dataArray_51_13_MPORT_mask) begin
      dataArray_51_13[dataArray_51_13_MPORT_addr] <= dataArray_51_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_14_MPORT_en & dataArray_51_14_MPORT_mask) begin
      dataArray_51_14[dataArray_51_14_MPORT_addr] <= dataArray_51_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_51_15_MPORT_en & dataArray_51_15_MPORT_mask) begin
      dataArray_51_15[dataArray_51_15_MPORT_addr] <= dataArray_51_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_51_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_51_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_51_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_51_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_0_MPORT_en & dataArray_52_0_MPORT_mask) begin
      dataArray_52_0[dataArray_52_0_MPORT_addr] <= dataArray_52_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_1_MPORT_en & dataArray_52_1_MPORT_mask) begin
      dataArray_52_1[dataArray_52_1_MPORT_addr] <= dataArray_52_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_2_MPORT_en & dataArray_52_2_MPORT_mask) begin
      dataArray_52_2[dataArray_52_2_MPORT_addr] <= dataArray_52_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_3_MPORT_en & dataArray_52_3_MPORT_mask) begin
      dataArray_52_3[dataArray_52_3_MPORT_addr] <= dataArray_52_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_4_MPORT_en & dataArray_52_4_MPORT_mask) begin
      dataArray_52_4[dataArray_52_4_MPORT_addr] <= dataArray_52_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_5_MPORT_en & dataArray_52_5_MPORT_mask) begin
      dataArray_52_5[dataArray_52_5_MPORT_addr] <= dataArray_52_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_6_MPORT_en & dataArray_52_6_MPORT_mask) begin
      dataArray_52_6[dataArray_52_6_MPORT_addr] <= dataArray_52_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_7_MPORT_en & dataArray_52_7_MPORT_mask) begin
      dataArray_52_7[dataArray_52_7_MPORT_addr] <= dataArray_52_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_8_MPORT_en & dataArray_52_8_MPORT_mask) begin
      dataArray_52_8[dataArray_52_8_MPORT_addr] <= dataArray_52_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_9_MPORT_en & dataArray_52_9_MPORT_mask) begin
      dataArray_52_9[dataArray_52_9_MPORT_addr] <= dataArray_52_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_10_MPORT_en & dataArray_52_10_MPORT_mask) begin
      dataArray_52_10[dataArray_52_10_MPORT_addr] <= dataArray_52_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_11_MPORT_en & dataArray_52_11_MPORT_mask) begin
      dataArray_52_11[dataArray_52_11_MPORT_addr] <= dataArray_52_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_12_MPORT_en & dataArray_52_12_MPORT_mask) begin
      dataArray_52_12[dataArray_52_12_MPORT_addr] <= dataArray_52_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_13_MPORT_en & dataArray_52_13_MPORT_mask) begin
      dataArray_52_13[dataArray_52_13_MPORT_addr] <= dataArray_52_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_14_MPORT_en & dataArray_52_14_MPORT_mask) begin
      dataArray_52_14[dataArray_52_14_MPORT_addr] <= dataArray_52_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_52_15_MPORT_en & dataArray_52_15_MPORT_mask) begin
      dataArray_52_15[dataArray_52_15_MPORT_addr] <= dataArray_52_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_52_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_52_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_52_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_52_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_0_MPORT_en & dataArray_53_0_MPORT_mask) begin
      dataArray_53_0[dataArray_53_0_MPORT_addr] <= dataArray_53_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_1_MPORT_en & dataArray_53_1_MPORT_mask) begin
      dataArray_53_1[dataArray_53_1_MPORT_addr] <= dataArray_53_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_2_MPORT_en & dataArray_53_2_MPORT_mask) begin
      dataArray_53_2[dataArray_53_2_MPORT_addr] <= dataArray_53_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_3_MPORT_en & dataArray_53_3_MPORT_mask) begin
      dataArray_53_3[dataArray_53_3_MPORT_addr] <= dataArray_53_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_4_MPORT_en & dataArray_53_4_MPORT_mask) begin
      dataArray_53_4[dataArray_53_4_MPORT_addr] <= dataArray_53_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_5_MPORT_en & dataArray_53_5_MPORT_mask) begin
      dataArray_53_5[dataArray_53_5_MPORT_addr] <= dataArray_53_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_6_MPORT_en & dataArray_53_6_MPORT_mask) begin
      dataArray_53_6[dataArray_53_6_MPORT_addr] <= dataArray_53_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_7_MPORT_en & dataArray_53_7_MPORT_mask) begin
      dataArray_53_7[dataArray_53_7_MPORT_addr] <= dataArray_53_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_8_MPORT_en & dataArray_53_8_MPORT_mask) begin
      dataArray_53_8[dataArray_53_8_MPORT_addr] <= dataArray_53_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_9_MPORT_en & dataArray_53_9_MPORT_mask) begin
      dataArray_53_9[dataArray_53_9_MPORT_addr] <= dataArray_53_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_10_MPORT_en & dataArray_53_10_MPORT_mask) begin
      dataArray_53_10[dataArray_53_10_MPORT_addr] <= dataArray_53_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_11_MPORT_en & dataArray_53_11_MPORT_mask) begin
      dataArray_53_11[dataArray_53_11_MPORT_addr] <= dataArray_53_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_12_MPORT_en & dataArray_53_12_MPORT_mask) begin
      dataArray_53_12[dataArray_53_12_MPORT_addr] <= dataArray_53_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_13_MPORT_en & dataArray_53_13_MPORT_mask) begin
      dataArray_53_13[dataArray_53_13_MPORT_addr] <= dataArray_53_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_14_MPORT_en & dataArray_53_14_MPORT_mask) begin
      dataArray_53_14[dataArray_53_14_MPORT_addr] <= dataArray_53_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_53_15_MPORT_en & dataArray_53_15_MPORT_mask) begin
      dataArray_53_15[dataArray_53_15_MPORT_addr] <= dataArray_53_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_53_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_53_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_53_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_53_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_0_MPORT_en & dataArray_54_0_MPORT_mask) begin
      dataArray_54_0[dataArray_54_0_MPORT_addr] <= dataArray_54_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_1_MPORT_en & dataArray_54_1_MPORT_mask) begin
      dataArray_54_1[dataArray_54_1_MPORT_addr] <= dataArray_54_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_2_MPORT_en & dataArray_54_2_MPORT_mask) begin
      dataArray_54_2[dataArray_54_2_MPORT_addr] <= dataArray_54_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_3_MPORT_en & dataArray_54_3_MPORT_mask) begin
      dataArray_54_3[dataArray_54_3_MPORT_addr] <= dataArray_54_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_4_MPORT_en & dataArray_54_4_MPORT_mask) begin
      dataArray_54_4[dataArray_54_4_MPORT_addr] <= dataArray_54_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_5_MPORT_en & dataArray_54_5_MPORT_mask) begin
      dataArray_54_5[dataArray_54_5_MPORT_addr] <= dataArray_54_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_6_MPORT_en & dataArray_54_6_MPORT_mask) begin
      dataArray_54_6[dataArray_54_6_MPORT_addr] <= dataArray_54_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_7_MPORT_en & dataArray_54_7_MPORT_mask) begin
      dataArray_54_7[dataArray_54_7_MPORT_addr] <= dataArray_54_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_8_MPORT_en & dataArray_54_8_MPORT_mask) begin
      dataArray_54_8[dataArray_54_8_MPORT_addr] <= dataArray_54_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_9_MPORT_en & dataArray_54_9_MPORT_mask) begin
      dataArray_54_9[dataArray_54_9_MPORT_addr] <= dataArray_54_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_10_MPORT_en & dataArray_54_10_MPORT_mask) begin
      dataArray_54_10[dataArray_54_10_MPORT_addr] <= dataArray_54_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_11_MPORT_en & dataArray_54_11_MPORT_mask) begin
      dataArray_54_11[dataArray_54_11_MPORT_addr] <= dataArray_54_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_12_MPORT_en & dataArray_54_12_MPORT_mask) begin
      dataArray_54_12[dataArray_54_12_MPORT_addr] <= dataArray_54_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_13_MPORT_en & dataArray_54_13_MPORT_mask) begin
      dataArray_54_13[dataArray_54_13_MPORT_addr] <= dataArray_54_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_14_MPORT_en & dataArray_54_14_MPORT_mask) begin
      dataArray_54_14[dataArray_54_14_MPORT_addr] <= dataArray_54_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_54_15_MPORT_en & dataArray_54_15_MPORT_mask) begin
      dataArray_54_15[dataArray_54_15_MPORT_addr] <= dataArray_54_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_54_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_54_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_54_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_54_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_0_MPORT_en & dataArray_55_0_MPORT_mask) begin
      dataArray_55_0[dataArray_55_0_MPORT_addr] <= dataArray_55_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_1_MPORT_en & dataArray_55_1_MPORT_mask) begin
      dataArray_55_1[dataArray_55_1_MPORT_addr] <= dataArray_55_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_2_MPORT_en & dataArray_55_2_MPORT_mask) begin
      dataArray_55_2[dataArray_55_2_MPORT_addr] <= dataArray_55_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_3_MPORT_en & dataArray_55_3_MPORT_mask) begin
      dataArray_55_3[dataArray_55_3_MPORT_addr] <= dataArray_55_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_4_MPORT_en & dataArray_55_4_MPORT_mask) begin
      dataArray_55_4[dataArray_55_4_MPORT_addr] <= dataArray_55_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_5_MPORT_en & dataArray_55_5_MPORT_mask) begin
      dataArray_55_5[dataArray_55_5_MPORT_addr] <= dataArray_55_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_6_MPORT_en & dataArray_55_6_MPORT_mask) begin
      dataArray_55_6[dataArray_55_6_MPORT_addr] <= dataArray_55_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_7_MPORT_en & dataArray_55_7_MPORT_mask) begin
      dataArray_55_7[dataArray_55_7_MPORT_addr] <= dataArray_55_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_8_MPORT_en & dataArray_55_8_MPORT_mask) begin
      dataArray_55_8[dataArray_55_8_MPORT_addr] <= dataArray_55_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_9_MPORT_en & dataArray_55_9_MPORT_mask) begin
      dataArray_55_9[dataArray_55_9_MPORT_addr] <= dataArray_55_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_10_MPORT_en & dataArray_55_10_MPORT_mask) begin
      dataArray_55_10[dataArray_55_10_MPORT_addr] <= dataArray_55_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_11_MPORT_en & dataArray_55_11_MPORT_mask) begin
      dataArray_55_11[dataArray_55_11_MPORT_addr] <= dataArray_55_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_12_MPORT_en & dataArray_55_12_MPORT_mask) begin
      dataArray_55_12[dataArray_55_12_MPORT_addr] <= dataArray_55_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_13_MPORT_en & dataArray_55_13_MPORT_mask) begin
      dataArray_55_13[dataArray_55_13_MPORT_addr] <= dataArray_55_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_14_MPORT_en & dataArray_55_14_MPORT_mask) begin
      dataArray_55_14[dataArray_55_14_MPORT_addr] <= dataArray_55_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_55_15_MPORT_en & dataArray_55_15_MPORT_mask) begin
      dataArray_55_15[dataArray_55_15_MPORT_addr] <= dataArray_55_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_55_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_55_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_55_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_55_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_0_MPORT_en & dataArray_56_0_MPORT_mask) begin
      dataArray_56_0[dataArray_56_0_MPORT_addr] <= dataArray_56_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_1_MPORT_en & dataArray_56_1_MPORT_mask) begin
      dataArray_56_1[dataArray_56_1_MPORT_addr] <= dataArray_56_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_2_MPORT_en & dataArray_56_2_MPORT_mask) begin
      dataArray_56_2[dataArray_56_2_MPORT_addr] <= dataArray_56_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_3_MPORT_en & dataArray_56_3_MPORT_mask) begin
      dataArray_56_3[dataArray_56_3_MPORT_addr] <= dataArray_56_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_4_MPORT_en & dataArray_56_4_MPORT_mask) begin
      dataArray_56_4[dataArray_56_4_MPORT_addr] <= dataArray_56_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_5_MPORT_en & dataArray_56_5_MPORT_mask) begin
      dataArray_56_5[dataArray_56_5_MPORT_addr] <= dataArray_56_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_6_MPORT_en & dataArray_56_6_MPORT_mask) begin
      dataArray_56_6[dataArray_56_6_MPORT_addr] <= dataArray_56_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_7_MPORT_en & dataArray_56_7_MPORT_mask) begin
      dataArray_56_7[dataArray_56_7_MPORT_addr] <= dataArray_56_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_8_MPORT_en & dataArray_56_8_MPORT_mask) begin
      dataArray_56_8[dataArray_56_8_MPORT_addr] <= dataArray_56_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_9_MPORT_en & dataArray_56_9_MPORT_mask) begin
      dataArray_56_9[dataArray_56_9_MPORT_addr] <= dataArray_56_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_10_MPORT_en & dataArray_56_10_MPORT_mask) begin
      dataArray_56_10[dataArray_56_10_MPORT_addr] <= dataArray_56_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_11_MPORT_en & dataArray_56_11_MPORT_mask) begin
      dataArray_56_11[dataArray_56_11_MPORT_addr] <= dataArray_56_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_12_MPORT_en & dataArray_56_12_MPORT_mask) begin
      dataArray_56_12[dataArray_56_12_MPORT_addr] <= dataArray_56_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_13_MPORT_en & dataArray_56_13_MPORT_mask) begin
      dataArray_56_13[dataArray_56_13_MPORT_addr] <= dataArray_56_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_14_MPORT_en & dataArray_56_14_MPORT_mask) begin
      dataArray_56_14[dataArray_56_14_MPORT_addr] <= dataArray_56_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_56_15_MPORT_en & dataArray_56_15_MPORT_mask) begin
      dataArray_56_15[dataArray_56_15_MPORT_addr] <= dataArray_56_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_56_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_56_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_56_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_56_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_0_MPORT_en & dataArray_57_0_MPORT_mask) begin
      dataArray_57_0[dataArray_57_0_MPORT_addr] <= dataArray_57_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_1_MPORT_en & dataArray_57_1_MPORT_mask) begin
      dataArray_57_1[dataArray_57_1_MPORT_addr] <= dataArray_57_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_2_MPORT_en & dataArray_57_2_MPORT_mask) begin
      dataArray_57_2[dataArray_57_2_MPORT_addr] <= dataArray_57_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_3_MPORT_en & dataArray_57_3_MPORT_mask) begin
      dataArray_57_3[dataArray_57_3_MPORT_addr] <= dataArray_57_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_4_MPORT_en & dataArray_57_4_MPORT_mask) begin
      dataArray_57_4[dataArray_57_4_MPORT_addr] <= dataArray_57_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_5_MPORT_en & dataArray_57_5_MPORT_mask) begin
      dataArray_57_5[dataArray_57_5_MPORT_addr] <= dataArray_57_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_6_MPORT_en & dataArray_57_6_MPORT_mask) begin
      dataArray_57_6[dataArray_57_6_MPORT_addr] <= dataArray_57_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_7_MPORT_en & dataArray_57_7_MPORT_mask) begin
      dataArray_57_7[dataArray_57_7_MPORT_addr] <= dataArray_57_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_8_MPORT_en & dataArray_57_8_MPORT_mask) begin
      dataArray_57_8[dataArray_57_8_MPORT_addr] <= dataArray_57_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_9_MPORT_en & dataArray_57_9_MPORT_mask) begin
      dataArray_57_9[dataArray_57_9_MPORT_addr] <= dataArray_57_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_10_MPORT_en & dataArray_57_10_MPORT_mask) begin
      dataArray_57_10[dataArray_57_10_MPORT_addr] <= dataArray_57_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_11_MPORT_en & dataArray_57_11_MPORT_mask) begin
      dataArray_57_11[dataArray_57_11_MPORT_addr] <= dataArray_57_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_12_MPORT_en & dataArray_57_12_MPORT_mask) begin
      dataArray_57_12[dataArray_57_12_MPORT_addr] <= dataArray_57_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_13_MPORT_en & dataArray_57_13_MPORT_mask) begin
      dataArray_57_13[dataArray_57_13_MPORT_addr] <= dataArray_57_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_14_MPORT_en & dataArray_57_14_MPORT_mask) begin
      dataArray_57_14[dataArray_57_14_MPORT_addr] <= dataArray_57_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_57_15_MPORT_en & dataArray_57_15_MPORT_mask) begin
      dataArray_57_15[dataArray_57_15_MPORT_addr] <= dataArray_57_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_57_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_57_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_57_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_57_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_0_MPORT_en & dataArray_58_0_MPORT_mask) begin
      dataArray_58_0[dataArray_58_0_MPORT_addr] <= dataArray_58_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_1_MPORT_en & dataArray_58_1_MPORT_mask) begin
      dataArray_58_1[dataArray_58_1_MPORT_addr] <= dataArray_58_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_2_MPORT_en & dataArray_58_2_MPORT_mask) begin
      dataArray_58_2[dataArray_58_2_MPORT_addr] <= dataArray_58_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_3_MPORT_en & dataArray_58_3_MPORT_mask) begin
      dataArray_58_3[dataArray_58_3_MPORT_addr] <= dataArray_58_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_4_MPORT_en & dataArray_58_4_MPORT_mask) begin
      dataArray_58_4[dataArray_58_4_MPORT_addr] <= dataArray_58_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_5_MPORT_en & dataArray_58_5_MPORT_mask) begin
      dataArray_58_5[dataArray_58_5_MPORT_addr] <= dataArray_58_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_6_MPORT_en & dataArray_58_6_MPORT_mask) begin
      dataArray_58_6[dataArray_58_6_MPORT_addr] <= dataArray_58_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_7_MPORT_en & dataArray_58_7_MPORT_mask) begin
      dataArray_58_7[dataArray_58_7_MPORT_addr] <= dataArray_58_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_8_MPORT_en & dataArray_58_8_MPORT_mask) begin
      dataArray_58_8[dataArray_58_8_MPORT_addr] <= dataArray_58_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_9_MPORT_en & dataArray_58_9_MPORT_mask) begin
      dataArray_58_9[dataArray_58_9_MPORT_addr] <= dataArray_58_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_10_MPORT_en & dataArray_58_10_MPORT_mask) begin
      dataArray_58_10[dataArray_58_10_MPORT_addr] <= dataArray_58_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_11_MPORT_en & dataArray_58_11_MPORT_mask) begin
      dataArray_58_11[dataArray_58_11_MPORT_addr] <= dataArray_58_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_12_MPORT_en & dataArray_58_12_MPORT_mask) begin
      dataArray_58_12[dataArray_58_12_MPORT_addr] <= dataArray_58_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_13_MPORT_en & dataArray_58_13_MPORT_mask) begin
      dataArray_58_13[dataArray_58_13_MPORT_addr] <= dataArray_58_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_14_MPORT_en & dataArray_58_14_MPORT_mask) begin
      dataArray_58_14[dataArray_58_14_MPORT_addr] <= dataArray_58_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_58_15_MPORT_en & dataArray_58_15_MPORT_mask) begin
      dataArray_58_15[dataArray_58_15_MPORT_addr] <= dataArray_58_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_58_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_58_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_58_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_58_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_0_MPORT_en & dataArray_59_0_MPORT_mask) begin
      dataArray_59_0[dataArray_59_0_MPORT_addr] <= dataArray_59_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_1_MPORT_en & dataArray_59_1_MPORT_mask) begin
      dataArray_59_1[dataArray_59_1_MPORT_addr] <= dataArray_59_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_2_MPORT_en & dataArray_59_2_MPORT_mask) begin
      dataArray_59_2[dataArray_59_2_MPORT_addr] <= dataArray_59_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_3_MPORT_en & dataArray_59_3_MPORT_mask) begin
      dataArray_59_3[dataArray_59_3_MPORT_addr] <= dataArray_59_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_4_MPORT_en & dataArray_59_4_MPORT_mask) begin
      dataArray_59_4[dataArray_59_4_MPORT_addr] <= dataArray_59_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_5_MPORT_en & dataArray_59_5_MPORT_mask) begin
      dataArray_59_5[dataArray_59_5_MPORT_addr] <= dataArray_59_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_6_MPORT_en & dataArray_59_6_MPORT_mask) begin
      dataArray_59_6[dataArray_59_6_MPORT_addr] <= dataArray_59_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_7_MPORT_en & dataArray_59_7_MPORT_mask) begin
      dataArray_59_7[dataArray_59_7_MPORT_addr] <= dataArray_59_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_8_MPORT_en & dataArray_59_8_MPORT_mask) begin
      dataArray_59_8[dataArray_59_8_MPORT_addr] <= dataArray_59_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_9_MPORT_en & dataArray_59_9_MPORT_mask) begin
      dataArray_59_9[dataArray_59_9_MPORT_addr] <= dataArray_59_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_10_MPORT_en & dataArray_59_10_MPORT_mask) begin
      dataArray_59_10[dataArray_59_10_MPORT_addr] <= dataArray_59_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_11_MPORT_en & dataArray_59_11_MPORT_mask) begin
      dataArray_59_11[dataArray_59_11_MPORT_addr] <= dataArray_59_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_12_MPORT_en & dataArray_59_12_MPORT_mask) begin
      dataArray_59_12[dataArray_59_12_MPORT_addr] <= dataArray_59_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_13_MPORT_en & dataArray_59_13_MPORT_mask) begin
      dataArray_59_13[dataArray_59_13_MPORT_addr] <= dataArray_59_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_14_MPORT_en & dataArray_59_14_MPORT_mask) begin
      dataArray_59_14[dataArray_59_14_MPORT_addr] <= dataArray_59_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_59_15_MPORT_en & dataArray_59_15_MPORT_mask) begin
      dataArray_59_15[dataArray_59_15_MPORT_addr] <= dataArray_59_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_59_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_59_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_59_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_59_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_0_MPORT_en & dataArray_60_0_MPORT_mask) begin
      dataArray_60_0[dataArray_60_0_MPORT_addr] <= dataArray_60_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_1_MPORT_en & dataArray_60_1_MPORT_mask) begin
      dataArray_60_1[dataArray_60_1_MPORT_addr] <= dataArray_60_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_2_MPORT_en & dataArray_60_2_MPORT_mask) begin
      dataArray_60_2[dataArray_60_2_MPORT_addr] <= dataArray_60_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_3_MPORT_en & dataArray_60_3_MPORT_mask) begin
      dataArray_60_3[dataArray_60_3_MPORT_addr] <= dataArray_60_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_4_MPORT_en & dataArray_60_4_MPORT_mask) begin
      dataArray_60_4[dataArray_60_4_MPORT_addr] <= dataArray_60_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_5_MPORT_en & dataArray_60_5_MPORT_mask) begin
      dataArray_60_5[dataArray_60_5_MPORT_addr] <= dataArray_60_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_6_MPORT_en & dataArray_60_6_MPORT_mask) begin
      dataArray_60_6[dataArray_60_6_MPORT_addr] <= dataArray_60_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_7_MPORT_en & dataArray_60_7_MPORT_mask) begin
      dataArray_60_7[dataArray_60_7_MPORT_addr] <= dataArray_60_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_8_MPORT_en & dataArray_60_8_MPORT_mask) begin
      dataArray_60_8[dataArray_60_8_MPORT_addr] <= dataArray_60_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_9_MPORT_en & dataArray_60_9_MPORT_mask) begin
      dataArray_60_9[dataArray_60_9_MPORT_addr] <= dataArray_60_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_10_MPORT_en & dataArray_60_10_MPORT_mask) begin
      dataArray_60_10[dataArray_60_10_MPORT_addr] <= dataArray_60_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_11_MPORT_en & dataArray_60_11_MPORT_mask) begin
      dataArray_60_11[dataArray_60_11_MPORT_addr] <= dataArray_60_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_12_MPORT_en & dataArray_60_12_MPORT_mask) begin
      dataArray_60_12[dataArray_60_12_MPORT_addr] <= dataArray_60_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_13_MPORT_en & dataArray_60_13_MPORT_mask) begin
      dataArray_60_13[dataArray_60_13_MPORT_addr] <= dataArray_60_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_14_MPORT_en & dataArray_60_14_MPORT_mask) begin
      dataArray_60_14[dataArray_60_14_MPORT_addr] <= dataArray_60_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_60_15_MPORT_en & dataArray_60_15_MPORT_mask) begin
      dataArray_60_15[dataArray_60_15_MPORT_addr] <= dataArray_60_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_60_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_60_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_60_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_60_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_0_MPORT_en & dataArray_61_0_MPORT_mask) begin
      dataArray_61_0[dataArray_61_0_MPORT_addr] <= dataArray_61_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_1_MPORT_en & dataArray_61_1_MPORT_mask) begin
      dataArray_61_1[dataArray_61_1_MPORT_addr] <= dataArray_61_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_2_MPORT_en & dataArray_61_2_MPORT_mask) begin
      dataArray_61_2[dataArray_61_2_MPORT_addr] <= dataArray_61_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_3_MPORT_en & dataArray_61_3_MPORT_mask) begin
      dataArray_61_3[dataArray_61_3_MPORT_addr] <= dataArray_61_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_4_MPORT_en & dataArray_61_4_MPORT_mask) begin
      dataArray_61_4[dataArray_61_4_MPORT_addr] <= dataArray_61_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_5_MPORT_en & dataArray_61_5_MPORT_mask) begin
      dataArray_61_5[dataArray_61_5_MPORT_addr] <= dataArray_61_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_6_MPORT_en & dataArray_61_6_MPORT_mask) begin
      dataArray_61_6[dataArray_61_6_MPORT_addr] <= dataArray_61_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_7_MPORT_en & dataArray_61_7_MPORT_mask) begin
      dataArray_61_7[dataArray_61_7_MPORT_addr] <= dataArray_61_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_8_MPORT_en & dataArray_61_8_MPORT_mask) begin
      dataArray_61_8[dataArray_61_8_MPORT_addr] <= dataArray_61_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_9_MPORT_en & dataArray_61_9_MPORT_mask) begin
      dataArray_61_9[dataArray_61_9_MPORT_addr] <= dataArray_61_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_10_MPORT_en & dataArray_61_10_MPORT_mask) begin
      dataArray_61_10[dataArray_61_10_MPORT_addr] <= dataArray_61_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_11_MPORT_en & dataArray_61_11_MPORT_mask) begin
      dataArray_61_11[dataArray_61_11_MPORT_addr] <= dataArray_61_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_12_MPORT_en & dataArray_61_12_MPORT_mask) begin
      dataArray_61_12[dataArray_61_12_MPORT_addr] <= dataArray_61_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_13_MPORT_en & dataArray_61_13_MPORT_mask) begin
      dataArray_61_13[dataArray_61_13_MPORT_addr] <= dataArray_61_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_14_MPORT_en & dataArray_61_14_MPORT_mask) begin
      dataArray_61_14[dataArray_61_14_MPORT_addr] <= dataArray_61_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_61_15_MPORT_en & dataArray_61_15_MPORT_mask) begin
      dataArray_61_15[dataArray_61_15_MPORT_addr] <= dataArray_61_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_61_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_61_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_61_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_61_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_0_MPORT_en & dataArray_62_0_MPORT_mask) begin
      dataArray_62_0[dataArray_62_0_MPORT_addr] <= dataArray_62_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_1_MPORT_en & dataArray_62_1_MPORT_mask) begin
      dataArray_62_1[dataArray_62_1_MPORT_addr] <= dataArray_62_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_2_MPORT_en & dataArray_62_2_MPORT_mask) begin
      dataArray_62_2[dataArray_62_2_MPORT_addr] <= dataArray_62_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_3_MPORT_en & dataArray_62_3_MPORT_mask) begin
      dataArray_62_3[dataArray_62_3_MPORT_addr] <= dataArray_62_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_4_MPORT_en & dataArray_62_4_MPORT_mask) begin
      dataArray_62_4[dataArray_62_4_MPORT_addr] <= dataArray_62_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_5_MPORT_en & dataArray_62_5_MPORT_mask) begin
      dataArray_62_5[dataArray_62_5_MPORT_addr] <= dataArray_62_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_6_MPORT_en & dataArray_62_6_MPORT_mask) begin
      dataArray_62_6[dataArray_62_6_MPORT_addr] <= dataArray_62_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_7_MPORT_en & dataArray_62_7_MPORT_mask) begin
      dataArray_62_7[dataArray_62_7_MPORT_addr] <= dataArray_62_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_8_MPORT_en & dataArray_62_8_MPORT_mask) begin
      dataArray_62_8[dataArray_62_8_MPORT_addr] <= dataArray_62_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_9_MPORT_en & dataArray_62_9_MPORT_mask) begin
      dataArray_62_9[dataArray_62_9_MPORT_addr] <= dataArray_62_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_10_MPORT_en & dataArray_62_10_MPORT_mask) begin
      dataArray_62_10[dataArray_62_10_MPORT_addr] <= dataArray_62_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_11_MPORT_en & dataArray_62_11_MPORT_mask) begin
      dataArray_62_11[dataArray_62_11_MPORT_addr] <= dataArray_62_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_12_MPORT_en & dataArray_62_12_MPORT_mask) begin
      dataArray_62_12[dataArray_62_12_MPORT_addr] <= dataArray_62_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_13_MPORT_en & dataArray_62_13_MPORT_mask) begin
      dataArray_62_13[dataArray_62_13_MPORT_addr] <= dataArray_62_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_14_MPORT_en & dataArray_62_14_MPORT_mask) begin
      dataArray_62_14[dataArray_62_14_MPORT_addr] <= dataArray_62_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_62_15_MPORT_en & dataArray_62_15_MPORT_mask) begin
      dataArray_62_15[dataArray_62_15_MPORT_addr] <= dataArray_62_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_62_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_62_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_62_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_62_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_0_MPORT_en & dataArray_63_0_MPORT_mask) begin
      dataArray_63_0[dataArray_63_0_MPORT_addr] <= dataArray_63_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_0_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_0_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_0_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_1_MPORT_en & dataArray_63_1_MPORT_mask) begin
      dataArray_63_1[dataArray_63_1_MPORT_addr] <= dataArray_63_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_1_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_1_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_1_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_2_MPORT_en & dataArray_63_2_MPORT_mask) begin
      dataArray_63_2[dataArray_63_2_MPORT_addr] <= dataArray_63_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_2_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_2_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_2_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_3_MPORT_en & dataArray_63_3_MPORT_mask) begin
      dataArray_63_3[dataArray_63_3_MPORT_addr] <= dataArray_63_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_3_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_3_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_3_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_4_MPORT_en & dataArray_63_4_MPORT_mask) begin
      dataArray_63_4[dataArray_63_4_MPORT_addr] <= dataArray_63_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_4_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_4_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_4_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_5_MPORT_en & dataArray_63_5_MPORT_mask) begin
      dataArray_63_5[dataArray_63_5_MPORT_addr] <= dataArray_63_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_5_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_5_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_5_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_6_MPORT_en & dataArray_63_6_MPORT_mask) begin
      dataArray_63_6[dataArray_63_6_MPORT_addr] <= dataArray_63_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_6_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_6_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_6_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_7_MPORT_en & dataArray_63_7_MPORT_mask) begin
      dataArray_63_7[dataArray_63_7_MPORT_addr] <= dataArray_63_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_7_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_7_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_7_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_8_MPORT_en & dataArray_63_8_MPORT_mask) begin
      dataArray_63_8[dataArray_63_8_MPORT_addr] <= dataArray_63_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_8_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_8_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_8_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_9_MPORT_en & dataArray_63_9_MPORT_mask) begin
      dataArray_63_9[dataArray_63_9_MPORT_addr] <= dataArray_63_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_9_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_9_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_9_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_10_MPORT_en & dataArray_63_10_MPORT_mask) begin
      dataArray_63_10[dataArray_63_10_MPORT_addr] <= dataArray_63_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_10_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_10_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_10_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_11_MPORT_en & dataArray_63_11_MPORT_mask) begin
      dataArray_63_11[dataArray_63_11_MPORT_addr] <= dataArray_63_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_11_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_11_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_11_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_12_MPORT_en & dataArray_63_12_MPORT_mask) begin
      dataArray_63_12[dataArray_63_12_MPORT_addr] <= dataArray_63_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_12_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_12_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_12_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_13_MPORT_en & dataArray_63_13_MPORT_mask) begin
      dataArray_63_13[dataArray_63_13_MPORT_addr] <= dataArray_63_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_13_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_13_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_13_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_14_MPORT_en & dataArray_63_14_MPORT_mask) begin
      dataArray_63_14[dataArray_63_14_MPORT_addr] <= dataArray_63_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_14_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_14_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_14_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (dataArray_63_15_MPORT_en & dataArray_63_15_MPORT_mask) begin
      dataArray_63_15[dataArray_63_15_MPORT_addr] <= dataArray_63_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_63_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (_SetId_T_6) begin
        dataArray_63_15_cachedata_MPORT_addr_pipe_0 <= 2'h3;
      end else if (_GEN_319 == tag) begin // @[Mux.scala 81:58]
        dataArray_63_15_cachedata_MPORT_addr_pipe_0 <= 2'h2;
      end else begin
        dataArray_63_15_cachedata_MPORT_addr_pipe_0 <= {{1'd0}, _GEN_191 == tag};
      end
    end
    if (reset) begin // @[cache.scala 21:30]
      replace_set <= 2'h0; // @[cache.scala 21:30]
    end else if (!(3'h0 == state_cache)) begin // @[cache.scala 49:26]
      if (!(3'h1 == state_cache)) begin // @[cache.scala 49:26]
        if (3'h2 == state_cache) begin // @[cache.scala 49:26]
          replace_set <= random_num; // @[cache.scala 64:25]
        end
      end
    end
    if (reset) begin // @[cache.scala 27:29]
      random_num <= 2'h0; // @[cache.scala 27:29]
    end else begin
      random_num <= _random_num_T_1; // @[cache.scala 28:16]
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_0 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7184) begin // @[cache.scala 84:50]
          tagArray_0_0 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_1 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7216) begin // @[cache.scala 84:50]
          tagArray_0_1 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_2 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7248) begin // @[cache.scala 84:50]
          tagArray_0_2 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_3 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7280) begin // @[cache.scala 84:50]
          tagArray_0_3 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_4 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7312) begin // @[cache.scala 84:50]
          tagArray_0_4 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_5 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7344) begin // @[cache.scala 84:50]
          tagArray_0_5 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_6 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7376) begin // @[cache.scala 84:50]
          tagArray_0_6 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_7 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7408) begin // @[cache.scala 84:50]
          tagArray_0_7 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_8 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7440) begin // @[cache.scala 84:50]
          tagArray_0_8 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_9 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7472) begin // @[cache.scala 84:50]
          tagArray_0_9 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_10 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7504) begin // @[cache.scala 84:50]
          tagArray_0_10 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_11 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7536) begin // @[cache.scala 84:50]
          tagArray_0_11 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_12 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7568) begin // @[cache.scala 84:50]
          tagArray_0_12 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_13 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7600) begin // @[cache.scala 84:50]
          tagArray_0_13 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_14 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7632) begin // @[cache.scala 84:50]
          tagArray_0_14 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_15 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7664) begin // @[cache.scala 84:50]
          tagArray_0_15 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_16 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7696) begin // @[cache.scala 84:50]
          tagArray_0_16 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_17 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7728) begin // @[cache.scala 84:50]
          tagArray_0_17 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_18 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7760) begin // @[cache.scala 84:50]
          tagArray_0_18 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_19 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7792) begin // @[cache.scala 84:50]
          tagArray_0_19 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_20 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7824) begin // @[cache.scala 84:50]
          tagArray_0_20 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_21 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7856) begin // @[cache.scala 84:50]
          tagArray_0_21 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_22 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7888) begin // @[cache.scala 84:50]
          tagArray_0_22 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_23 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7920) begin // @[cache.scala 84:50]
          tagArray_0_23 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_24 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7952) begin // @[cache.scala 84:50]
          tagArray_0_24 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_25 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_7984) begin // @[cache.scala 84:50]
          tagArray_0_25 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_26 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8016) begin // @[cache.scala 84:50]
          tagArray_0_26 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_27 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8048) begin // @[cache.scala 84:50]
          tagArray_0_27 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_28 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8080) begin // @[cache.scala 84:50]
          tagArray_0_28 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_29 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8112) begin // @[cache.scala 84:50]
          tagArray_0_29 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_30 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8144) begin // @[cache.scala 84:50]
          tagArray_0_30 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_31 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8176) begin // @[cache.scala 84:50]
          tagArray_0_31 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_32 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8208) begin // @[cache.scala 84:50]
          tagArray_0_32 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_33 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8240) begin // @[cache.scala 84:50]
          tagArray_0_33 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_34 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8272) begin // @[cache.scala 84:50]
          tagArray_0_34 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_35 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8304) begin // @[cache.scala 84:50]
          tagArray_0_35 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_36 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8336) begin // @[cache.scala 84:50]
          tagArray_0_36 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_37 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8368) begin // @[cache.scala 84:50]
          tagArray_0_37 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_38 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8400) begin // @[cache.scala 84:50]
          tagArray_0_38 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_39 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8432) begin // @[cache.scala 84:50]
          tagArray_0_39 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_40 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8464) begin // @[cache.scala 84:50]
          tagArray_0_40 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_41 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8496) begin // @[cache.scala 84:50]
          tagArray_0_41 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_42 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8528) begin // @[cache.scala 84:50]
          tagArray_0_42 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_43 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8560) begin // @[cache.scala 84:50]
          tagArray_0_43 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_44 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8592) begin // @[cache.scala 84:50]
          tagArray_0_44 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_45 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8624) begin // @[cache.scala 84:50]
          tagArray_0_45 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_46 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8656) begin // @[cache.scala 84:50]
          tagArray_0_46 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_47 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8688) begin // @[cache.scala 84:50]
          tagArray_0_47 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_48 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8720) begin // @[cache.scala 84:50]
          tagArray_0_48 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_49 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8752) begin // @[cache.scala 84:50]
          tagArray_0_49 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_50 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8784) begin // @[cache.scala 84:50]
          tagArray_0_50 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_51 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8816) begin // @[cache.scala 84:50]
          tagArray_0_51 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_52 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8848) begin // @[cache.scala 84:50]
          tagArray_0_52 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_53 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8880) begin // @[cache.scala 84:50]
          tagArray_0_53 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_54 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8912) begin // @[cache.scala 84:50]
          tagArray_0_54 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_55 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8944) begin // @[cache.scala 84:50]
          tagArray_0_55 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_56 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_8976) begin // @[cache.scala 84:50]
          tagArray_0_56 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_57 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9008) begin // @[cache.scala 84:50]
          tagArray_0_57 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_58 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9040) begin // @[cache.scala 84:50]
          tagArray_0_58 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_59 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9072) begin // @[cache.scala 84:50]
          tagArray_0_59 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_60 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9104) begin // @[cache.scala 84:50]
          tagArray_0_60 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_61 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9136) begin // @[cache.scala 84:50]
          tagArray_0_61 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_62 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9168) begin // @[cache.scala 84:50]
          tagArray_0_62 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_63 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9232 & _GEN_9200) begin // @[cache.scala 84:50]
          tagArray_0_63 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_0 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7184) begin // @[cache.scala 84:50]
          tagArray_1_0 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_1 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7216) begin // @[cache.scala 84:50]
          tagArray_1_1 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_2 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7248) begin // @[cache.scala 84:50]
          tagArray_1_2 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_3 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7280) begin // @[cache.scala 84:50]
          tagArray_1_3 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_4 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7312) begin // @[cache.scala 84:50]
          tagArray_1_4 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_5 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7344) begin // @[cache.scala 84:50]
          tagArray_1_5 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_6 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7376) begin // @[cache.scala 84:50]
          tagArray_1_6 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_7 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7408) begin // @[cache.scala 84:50]
          tagArray_1_7 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_8 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7440) begin // @[cache.scala 84:50]
          tagArray_1_8 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_9 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7472) begin // @[cache.scala 84:50]
          tagArray_1_9 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_10 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7504) begin // @[cache.scala 84:50]
          tagArray_1_10 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_11 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7536) begin // @[cache.scala 84:50]
          tagArray_1_11 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_12 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7568) begin // @[cache.scala 84:50]
          tagArray_1_12 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_13 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7600) begin // @[cache.scala 84:50]
          tagArray_1_13 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_14 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7632) begin // @[cache.scala 84:50]
          tagArray_1_14 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_15 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7664) begin // @[cache.scala 84:50]
          tagArray_1_15 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_16 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7696) begin // @[cache.scala 84:50]
          tagArray_1_16 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_17 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7728) begin // @[cache.scala 84:50]
          tagArray_1_17 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_18 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7760) begin // @[cache.scala 84:50]
          tagArray_1_18 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_19 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7792) begin // @[cache.scala 84:50]
          tagArray_1_19 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_20 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7824) begin // @[cache.scala 84:50]
          tagArray_1_20 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_21 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7856) begin // @[cache.scala 84:50]
          tagArray_1_21 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_22 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7888) begin // @[cache.scala 84:50]
          tagArray_1_22 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_23 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7920) begin // @[cache.scala 84:50]
          tagArray_1_23 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_24 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7952) begin // @[cache.scala 84:50]
          tagArray_1_24 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_25 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_7984) begin // @[cache.scala 84:50]
          tagArray_1_25 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_26 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8016) begin // @[cache.scala 84:50]
          tagArray_1_26 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_27 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8048) begin // @[cache.scala 84:50]
          tagArray_1_27 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_28 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8080) begin // @[cache.scala 84:50]
          tagArray_1_28 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_29 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8112) begin // @[cache.scala 84:50]
          tagArray_1_29 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_30 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8144) begin // @[cache.scala 84:50]
          tagArray_1_30 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_31 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8176) begin // @[cache.scala 84:50]
          tagArray_1_31 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_32 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8208) begin // @[cache.scala 84:50]
          tagArray_1_32 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_33 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8240) begin // @[cache.scala 84:50]
          tagArray_1_33 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_34 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8272) begin // @[cache.scala 84:50]
          tagArray_1_34 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_35 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8304) begin // @[cache.scala 84:50]
          tagArray_1_35 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_36 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8336) begin // @[cache.scala 84:50]
          tagArray_1_36 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_37 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8368) begin // @[cache.scala 84:50]
          tagArray_1_37 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_38 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8400) begin // @[cache.scala 84:50]
          tagArray_1_38 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_39 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8432) begin // @[cache.scala 84:50]
          tagArray_1_39 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_40 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8464) begin // @[cache.scala 84:50]
          tagArray_1_40 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_41 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8496) begin // @[cache.scala 84:50]
          tagArray_1_41 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_42 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8528) begin // @[cache.scala 84:50]
          tagArray_1_42 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_43 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8560) begin // @[cache.scala 84:50]
          tagArray_1_43 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_44 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8592) begin // @[cache.scala 84:50]
          tagArray_1_44 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_45 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8624) begin // @[cache.scala 84:50]
          tagArray_1_45 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_46 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8656) begin // @[cache.scala 84:50]
          tagArray_1_46 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_47 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8688) begin // @[cache.scala 84:50]
          tagArray_1_47 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_48 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8720) begin // @[cache.scala 84:50]
          tagArray_1_48 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_49 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8752) begin // @[cache.scala 84:50]
          tagArray_1_49 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_50 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8784) begin // @[cache.scala 84:50]
          tagArray_1_50 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_51 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8816) begin // @[cache.scala 84:50]
          tagArray_1_51 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_52 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8848) begin // @[cache.scala 84:50]
          tagArray_1_52 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_53 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8880) begin // @[cache.scala 84:50]
          tagArray_1_53 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_54 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8912) begin // @[cache.scala 84:50]
          tagArray_1_54 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_55 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8944) begin // @[cache.scala 84:50]
          tagArray_1_55 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_56 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_8976) begin // @[cache.scala 84:50]
          tagArray_1_56 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_57 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9008) begin // @[cache.scala 84:50]
          tagArray_1_57 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_58 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9040) begin // @[cache.scala 84:50]
          tagArray_1_58 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_59 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9072) begin // @[cache.scala 84:50]
          tagArray_1_59 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_60 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9104) begin // @[cache.scala 84:50]
          tagArray_1_60 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_61 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9136) begin // @[cache.scala 84:50]
          tagArray_1_61 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_62 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9168) begin // @[cache.scala 84:50]
          tagArray_1_62 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_63 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9424 & _GEN_9200) begin // @[cache.scala 84:50]
          tagArray_1_63 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_0 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7184) begin // @[cache.scala 84:50]
          tagArray_2_0 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_1 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7216) begin // @[cache.scala 84:50]
          tagArray_2_1 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_2 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7248) begin // @[cache.scala 84:50]
          tagArray_2_2 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_3 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7280) begin // @[cache.scala 84:50]
          tagArray_2_3 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_4 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7312) begin // @[cache.scala 84:50]
          tagArray_2_4 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_5 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7344) begin // @[cache.scala 84:50]
          tagArray_2_5 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_6 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7376) begin // @[cache.scala 84:50]
          tagArray_2_6 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_7 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7408) begin // @[cache.scala 84:50]
          tagArray_2_7 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_8 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7440) begin // @[cache.scala 84:50]
          tagArray_2_8 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_9 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7472) begin // @[cache.scala 84:50]
          tagArray_2_9 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_10 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7504) begin // @[cache.scala 84:50]
          tagArray_2_10 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_11 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7536) begin // @[cache.scala 84:50]
          tagArray_2_11 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_12 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7568) begin // @[cache.scala 84:50]
          tagArray_2_12 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_13 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7600) begin // @[cache.scala 84:50]
          tagArray_2_13 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_14 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7632) begin // @[cache.scala 84:50]
          tagArray_2_14 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_15 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7664) begin // @[cache.scala 84:50]
          tagArray_2_15 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_16 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7696) begin // @[cache.scala 84:50]
          tagArray_2_16 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_17 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7728) begin // @[cache.scala 84:50]
          tagArray_2_17 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_18 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7760) begin // @[cache.scala 84:50]
          tagArray_2_18 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_19 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7792) begin // @[cache.scala 84:50]
          tagArray_2_19 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_20 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7824) begin // @[cache.scala 84:50]
          tagArray_2_20 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_21 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7856) begin // @[cache.scala 84:50]
          tagArray_2_21 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_22 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7888) begin // @[cache.scala 84:50]
          tagArray_2_22 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_23 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7920) begin // @[cache.scala 84:50]
          tagArray_2_23 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_24 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7952) begin // @[cache.scala 84:50]
          tagArray_2_24 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_25 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_7984) begin // @[cache.scala 84:50]
          tagArray_2_25 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_26 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8016) begin // @[cache.scala 84:50]
          tagArray_2_26 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_27 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8048) begin // @[cache.scala 84:50]
          tagArray_2_27 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_28 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8080) begin // @[cache.scala 84:50]
          tagArray_2_28 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_29 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8112) begin // @[cache.scala 84:50]
          tagArray_2_29 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_30 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8144) begin // @[cache.scala 84:50]
          tagArray_2_30 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_31 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8176) begin // @[cache.scala 84:50]
          tagArray_2_31 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_32 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8208) begin // @[cache.scala 84:50]
          tagArray_2_32 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_33 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8240) begin // @[cache.scala 84:50]
          tagArray_2_33 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_34 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8272) begin // @[cache.scala 84:50]
          tagArray_2_34 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_35 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8304) begin // @[cache.scala 84:50]
          tagArray_2_35 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_36 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8336) begin // @[cache.scala 84:50]
          tagArray_2_36 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_37 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8368) begin // @[cache.scala 84:50]
          tagArray_2_37 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_38 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8400) begin // @[cache.scala 84:50]
          tagArray_2_38 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_39 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8432) begin // @[cache.scala 84:50]
          tagArray_2_39 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_40 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8464) begin // @[cache.scala 84:50]
          tagArray_2_40 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_41 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8496) begin // @[cache.scala 84:50]
          tagArray_2_41 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_42 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8528) begin // @[cache.scala 84:50]
          tagArray_2_42 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_43 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8560) begin // @[cache.scala 84:50]
          tagArray_2_43 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_44 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8592) begin // @[cache.scala 84:50]
          tagArray_2_44 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_45 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8624) begin // @[cache.scala 84:50]
          tagArray_2_45 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_46 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8656) begin // @[cache.scala 84:50]
          tagArray_2_46 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_47 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8688) begin // @[cache.scala 84:50]
          tagArray_2_47 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_48 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8720) begin // @[cache.scala 84:50]
          tagArray_2_48 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_49 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8752) begin // @[cache.scala 84:50]
          tagArray_2_49 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_50 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8784) begin // @[cache.scala 84:50]
          tagArray_2_50 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_51 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8816) begin // @[cache.scala 84:50]
          tagArray_2_51 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_52 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8848) begin // @[cache.scala 84:50]
          tagArray_2_52 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_53 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8880) begin // @[cache.scala 84:50]
          tagArray_2_53 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_54 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8912) begin // @[cache.scala 84:50]
          tagArray_2_54 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_55 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8944) begin // @[cache.scala 84:50]
          tagArray_2_55 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_56 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_8976) begin // @[cache.scala 84:50]
          tagArray_2_56 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_57 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9008) begin // @[cache.scala 84:50]
          tagArray_2_57 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_58 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9040) begin // @[cache.scala 84:50]
          tagArray_2_58 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_59 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9072) begin // @[cache.scala 84:50]
          tagArray_2_59 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_60 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9104) begin // @[cache.scala 84:50]
          tagArray_2_60 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_61 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9136) begin // @[cache.scala 84:50]
          tagArray_2_61 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_62 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9168) begin // @[cache.scala 84:50]
          tagArray_2_62 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_2_63 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9616 & _GEN_9200) begin // @[cache.scala 84:50]
          tagArray_2_63 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_0 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7184) begin // @[cache.scala 84:50]
          tagArray_3_0 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_1 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7216) begin // @[cache.scala 84:50]
          tagArray_3_1 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_2 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7248) begin // @[cache.scala 84:50]
          tagArray_3_2 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_3 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7280) begin // @[cache.scala 84:50]
          tagArray_3_3 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_4 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7312) begin // @[cache.scala 84:50]
          tagArray_3_4 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_5 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7344) begin // @[cache.scala 84:50]
          tagArray_3_5 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_6 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7376) begin // @[cache.scala 84:50]
          tagArray_3_6 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_7 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7408) begin // @[cache.scala 84:50]
          tagArray_3_7 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_8 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7440) begin // @[cache.scala 84:50]
          tagArray_3_8 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_9 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7472) begin // @[cache.scala 84:50]
          tagArray_3_9 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_10 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7504) begin // @[cache.scala 84:50]
          tagArray_3_10 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_11 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7536) begin // @[cache.scala 84:50]
          tagArray_3_11 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_12 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7568) begin // @[cache.scala 84:50]
          tagArray_3_12 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_13 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7600) begin // @[cache.scala 84:50]
          tagArray_3_13 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_14 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7632) begin // @[cache.scala 84:50]
          tagArray_3_14 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_15 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7664) begin // @[cache.scala 84:50]
          tagArray_3_15 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_16 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7696) begin // @[cache.scala 84:50]
          tagArray_3_16 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_17 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7728) begin // @[cache.scala 84:50]
          tagArray_3_17 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_18 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7760) begin // @[cache.scala 84:50]
          tagArray_3_18 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_19 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7792) begin // @[cache.scala 84:50]
          tagArray_3_19 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_20 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7824) begin // @[cache.scala 84:50]
          tagArray_3_20 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_21 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7856) begin // @[cache.scala 84:50]
          tagArray_3_21 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_22 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7888) begin // @[cache.scala 84:50]
          tagArray_3_22 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_23 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7920) begin // @[cache.scala 84:50]
          tagArray_3_23 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_24 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7952) begin // @[cache.scala 84:50]
          tagArray_3_24 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_25 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_7984) begin // @[cache.scala 84:50]
          tagArray_3_25 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_26 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8016) begin // @[cache.scala 84:50]
          tagArray_3_26 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_27 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8048) begin // @[cache.scala 84:50]
          tagArray_3_27 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_28 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8080) begin // @[cache.scala 84:50]
          tagArray_3_28 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_29 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8112) begin // @[cache.scala 84:50]
          tagArray_3_29 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_30 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8144) begin // @[cache.scala 84:50]
          tagArray_3_30 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_31 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8176) begin // @[cache.scala 84:50]
          tagArray_3_31 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_32 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8208) begin // @[cache.scala 84:50]
          tagArray_3_32 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_33 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8240) begin // @[cache.scala 84:50]
          tagArray_3_33 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_34 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8272) begin // @[cache.scala 84:50]
          tagArray_3_34 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_35 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8304) begin // @[cache.scala 84:50]
          tagArray_3_35 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_36 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8336) begin // @[cache.scala 84:50]
          tagArray_3_36 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_37 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8368) begin // @[cache.scala 84:50]
          tagArray_3_37 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_38 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8400) begin // @[cache.scala 84:50]
          tagArray_3_38 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_39 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8432) begin // @[cache.scala 84:50]
          tagArray_3_39 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_40 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8464) begin // @[cache.scala 84:50]
          tagArray_3_40 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_41 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8496) begin // @[cache.scala 84:50]
          tagArray_3_41 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_42 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8528) begin // @[cache.scala 84:50]
          tagArray_3_42 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_43 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8560) begin // @[cache.scala 84:50]
          tagArray_3_43 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_44 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8592) begin // @[cache.scala 84:50]
          tagArray_3_44 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_45 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8624) begin // @[cache.scala 84:50]
          tagArray_3_45 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_46 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8656) begin // @[cache.scala 84:50]
          tagArray_3_46 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_47 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8688) begin // @[cache.scala 84:50]
          tagArray_3_47 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_48 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8720) begin // @[cache.scala 84:50]
          tagArray_3_48 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_49 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8752) begin // @[cache.scala 84:50]
          tagArray_3_49 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_50 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8784) begin // @[cache.scala 84:50]
          tagArray_3_50 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_51 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8816) begin // @[cache.scala 84:50]
          tagArray_3_51 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_52 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8848) begin // @[cache.scala 84:50]
          tagArray_3_52 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_53 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8880) begin // @[cache.scala 84:50]
          tagArray_3_53 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_54 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8912) begin // @[cache.scala 84:50]
          tagArray_3_54 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_55 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8944) begin // @[cache.scala 84:50]
          tagArray_3_55 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_56 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_8976) begin // @[cache.scala 84:50]
          tagArray_3_56 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_57 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9008) begin // @[cache.scala 84:50]
          tagArray_3_57 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_58 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9040) begin // @[cache.scala 84:50]
          tagArray_3_58 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_59 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9072) begin // @[cache.scala 84:50]
          tagArray_3_59 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_60 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9104) begin // @[cache.scala 84:50]
          tagArray_3_60 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_61 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9136) begin // @[cache.scala 84:50]
          tagArray_3_61 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_62 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9168) begin // @[cache.scala 84:50]
          tagArray_3_62 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_3_63 <= 20'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_9808 & _GEN_9200) begin // @[cache.scala 84:50]
          tagArray_3_63 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_0 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_0 <= _GEN_2573;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_1 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_1 <= _GEN_2574;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_2 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_2 <= _GEN_2575;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_3 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_3 <= _GEN_2576;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_4 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_4 <= _GEN_2577;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_5 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_5 <= _GEN_2578;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_6 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_6 <= _GEN_2579;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_7 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_7 <= _GEN_2580;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_8 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_8 <= _GEN_2581;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_9 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_9 <= _GEN_2582;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_10 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_10 <= _GEN_2583;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_11 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_11 <= _GEN_2584;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_12 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_12 <= _GEN_2585;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_13 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_13 <= _GEN_2586;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_14 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_14 <= _GEN_2587;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_15 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_15 <= _GEN_2588;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_16 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_16 <= _GEN_2589;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_17 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_17 <= _GEN_2590;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_18 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_18 <= _GEN_2591;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_19 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_19 <= _GEN_2592;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_20 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_20 <= _GEN_2593;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_21 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_21 <= _GEN_2594;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_22 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_22 <= _GEN_2595;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_23 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_23 <= _GEN_2596;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_24 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_24 <= _GEN_2597;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_25 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_25 <= _GEN_2598;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_26 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_26 <= _GEN_2599;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_27 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_27 <= _GEN_2600;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_28 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_28 <= _GEN_2601;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_29 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_29 <= _GEN_2602;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_30 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_30 <= _GEN_2603;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_31 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_31 <= _GEN_2604;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_32 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_32 <= _GEN_2605;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_33 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_33 <= _GEN_2606;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_34 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_34 <= _GEN_2607;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_35 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_35 <= _GEN_2608;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_36 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_36 <= _GEN_2609;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_37 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_37 <= _GEN_2610;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_38 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_38 <= _GEN_2611;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_39 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_39 <= _GEN_2612;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_40 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_40 <= _GEN_2613;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_41 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_41 <= _GEN_2614;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_42 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_42 <= _GEN_2615;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_43 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_43 <= _GEN_2616;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_44 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_44 <= _GEN_2617;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_45 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_45 <= _GEN_2618;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_46 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_46 <= _GEN_2619;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_47 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_47 <= _GEN_2620;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_48 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_48 <= _GEN_2621;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_49 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_49 <= _GEN_2622;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_50 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_50 <= _GEN_2623;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_51 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_51 <= _GEN_2624;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_52 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_52 <= _GEN_2625;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_53 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_53 <= _GEN_2626;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_54 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_54 <= _GEN_2627;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_55 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_55 <= _GEN_2628;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_56 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_56 <= _GEN_2629;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_57 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_57 <= _GEN_2630;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_58 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_58 <= _GEN_2631;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_59 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_59 <= _GEN_2632;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_60 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_60 <= _GEN_2633;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_61 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_61 <= _GEN_2634;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_62 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_62 <= _GEN_2635;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_63 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_63 <= _GEN_2636;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_0 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_0 <= _GEN_2637;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_1 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_1 <= _GEN_2638;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_2 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_2 <= _GEN_2639;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_3 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_3 <= _GEN_2640;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_4 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_4 <= _GEN_2641;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_5 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_5 <= _GEN_2642;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_6 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_6 <= _GEN_2643;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_7 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_7 <= _GEN_2644;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_8 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_8 <= _GEN_2645;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_9 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_9 <= _GEN_2646;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_10 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_10 <= _GEN_2647;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_11 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_11 <= _GEN_2648;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_12 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_12 <= _GEN_2649;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_13 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_13 <= _GEN_2650;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_14 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_14 <= _GEN_2651;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_15 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_15 <= _GEN_2652;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_16 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_16 <= _GEN_2653;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_17 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_17 <= _GEN_2654;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_18 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_18 <= _GEN_2655;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_19 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_19 <= _GEN_2656;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_20 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_20 <= _GEN_2657;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_21 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_21 <= _GEN_2658;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_22 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_22 <= _GEN_2659;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_23 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_23 <= _GEN_2660;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_24 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_24 <= _GEN_2661;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_25 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_25 <= _GEN_2662;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_26 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_26 <= _GEN_2663;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_27 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_27 <= _GEN_2664;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_28 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_28 <= _GEN_2665;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_29 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_29 <= _GEN_2666;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_30 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_30 <= _GEN_2667;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_31 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_31 <= _GEN_2668;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_32 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_32 <= _GEN_2669;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_33 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_33 <= _GEN_2670;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_34 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_34 <= _GEN_2671;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_35 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_35 <= _GEN_2672;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_36 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_36 <= _GEN_2673;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_37 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_37 <= _GEN_2674;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_38 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_38 <= _GEN_2675;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_39 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_39 <= _GEN_2676;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_40 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_40 <= _GEN_2677;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_41 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_41 <= _GEN_2678;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_42 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_42 <= _GEN_2679;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_43 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_43 <= _GEN_2680;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_44 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_44 <= _GEN_2681;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_45 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_45 <= _GEN_2682;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_46 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_46 <= _GEN_2683;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_47 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_47 <= _GEN_2684;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_48 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_48 <= _GEN_2685;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_49 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_49 <= _GEN_2686;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_50 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_50 <= _GEN_2687;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_51 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_51 <= _GEN_2688;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_52 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_52 <= _GEN_2689;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_53 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_53 <= _GEN_2690;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_54 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_54 <= _GEN_2691;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_55 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_55 <= _GEN_2692;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_56 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_56 <= _GEN_2693;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_57 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_57 <= _GEN_2694;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_58 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_58 <= _GEN_2695;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_59 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_59 <= _GEN_2696;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_60 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_60 <= _GEN_2697;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_61 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_61 <= _GEN_2698;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_62 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_62 <= _GEN_2699;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_63 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_63 <= _GEN_2700;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_0 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_0 <= _GEN_2701;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_1 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_1 <= _GEN_2702;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_2 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_2 <= _GEN_2703;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_3 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_3 <= _GEN_2704;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_4 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_4 <= _GEN_2705;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_5 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_5 <= _GEN_2706;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_6 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_6 <= _GEN_2707;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_7 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_7 <= _GEN_2708;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_8 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_8 <= _GEN_2709;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_9 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_9 <= _GEN_2710;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_10 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_10 <= _GEN_2711;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_11 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_11 <= _GEN_2712;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_12 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_12 <= _GEN_2713;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_13 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_13 <= _GEN_2714;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_14 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_14 <= _GEN_2715;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_15 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_15 <= _GEN_2716;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_16 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_16 <= _GEN_2717;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_17 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_17 <= _GEN_2718;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_18 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_18 <= _GEN_2719;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_19 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_19 <= _GEN_2720;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_20 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_20 <= _GEN_2721;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_21 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_21 <= _GEN_2722;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_22 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_22 <= _GEN_2723;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_23 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_23 <= _GEN_2724;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_24 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_24 <= _GEN_2725;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_25 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_25 <= _GEN_2726;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_26 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_26 <= _GEN_2727;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_27 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_27 <= _GEN_2728;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_28 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_28 <= _GEN_2729;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_29 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_29 <= _GEN_2730;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_30 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_30 <= _GEN_2731;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_31 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_31 <= _GEN_2732;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_32 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_32 <= _GEN_2733;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_33 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_33 <= _GEN_2734;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_34 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_34 <= _GEN_2735;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_35 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_35 <= _GEN_2736;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_36 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_36 <= _GEN_2737;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_37 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_37 <= _GEN_2738;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_38 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_38 <= _GEN_2739;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_39 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_39 <= _GEN_2740;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_40 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_40 <= _GEN_2741;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_41 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_41 <= _GEN_2742;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_42 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_42 <= _GEN_2743;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_43 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_43 <= _GEN_2744;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_44 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_44 <= _GEN_2745;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_45 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_45 <= _GEN_2746;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_46 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_46 <= _GEN_2747;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_47 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_47 <= _GEN_2748;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_48 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_48 <= _GEN_2749;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_49 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_49 <= _GEN_2750;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_50 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_50 <= _GEN_2751;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_51 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_51 <= _GEN_2752;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_52 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_52 <= _GEN_2753;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_53 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_53 <= _GEN_2754;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_54 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_54 <= _GEN_2755;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_55 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_55 <= _GEN_2756;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_56 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_56 <= _GEN_2757;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_57 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_57 <= _GEN_2758;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_58 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_58 <= _GEN_2759;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_59 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_59 <= _GEN_2760;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_60 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_60 <= _GEN_2761;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_61 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_61 <= _GEN_2762;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_62 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_62 <= _GEN_2763;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_2_63 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_2_63 <= _GEN_2764;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_0 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_0 <= _GEN_2765;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_1 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_1 <= _GEN_2766;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_2 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_2 <= _GEN_2767;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_3 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_3 <= _GEN_2768;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_4 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_4 <= _GEN_2769;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_5 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_5 <= _GEN_2770;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_6 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_6 <= _GEN_2771;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_7 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_7 <= _GEN_2772;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_8 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_8 <= _GEN_2773;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_9 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_9 <= _GEN_2774;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_10 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_10 <= _GEN_2775;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_11 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_11 <= _GEN_2776;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_12 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_12 <= _GEN_2777;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_13 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_13 <= _GEN_2778;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_14 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_14 <= _GEN_2779;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_15 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_15 <= _GEN_2780;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_16 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_16 <= _GEN_2781;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_17 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_17 <= _GEN_2782;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_18 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_18 <= _GEN_2783;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_19 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_19 <= _GEN_2784;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_20 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_20 <= _GEN_2785;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_21 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_21 <= _GEN_2786;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_22 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_22 <= _GEN_2787;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_23 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_23 <= _GEN_2788;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_24 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_24 <= _GEN_2789;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_25 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_25 <= _GEN_2790;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_26 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_26 <= _GEN_2791;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_27 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_27 <= _GEN_2792;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_28 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_28 <= _GEN_2793;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_29 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_29 <= _GEN_2794;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_30 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_30 <= _GEN_2795;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_31 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_31 <= _GEN_2796;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_32 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_32 <= _GEN_2797;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_33 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_33 <= _GEN_2798;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_34 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_34 <= _GEN_2799;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_35 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_35 <= _GEN_2800;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_36 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_36 <= _GEN_2801;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_37 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_37 <= _GEN_2802;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_38 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_38 <= _GEN_2803;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_39 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_39 <= _GEN_2804;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_40 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_40 <= _GEN_2805;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_41 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_41 <= _GEN_2806;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_42 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_42 <= _GEN_2807;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_43 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_43 <= _GEN_2808;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_44 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_44 <= _GEN_2809;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_45 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_45 <= _GEN_2810;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_46 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_46 <= _GEN_2811;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_47 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_47 <= _GEN_2812;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_48 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_48 <= _GEN_2813;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_49 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_49 <= _GEN_2814;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_50 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_50 <= _GEN_2815;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_51 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_51 <= _GEN_2816;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_52 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_52 <= _GEN_2817;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_53 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_53 <= _GEN_2818;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_54 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_54 <= _GEN_2819;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_55 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_55 <= _GEN_2820;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_56 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_56 <= _GEN_2821;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_57 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_57 <= _GEN_2822;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_58 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_58 <= _GEN_2823;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_59 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_59 <= _GEN_2824;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_60 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_60 <= _GEN_2825;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_61 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_61 <= _GEN_2826;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_62 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_62 <= _GEN_2827;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_3_63 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_3_63 <= _GEN_2828;
      end
    end
    if (reset) begin // @[cache.scala 45:24]
      off <= 4'h0; // @[cache.scala 45:24]
    end else if (!(3'h0 == state_cache)) begin // @[cache.scala 49:26]
      if (!(3'h1 == state_cache)) begin // @[cache.scala 49:26]
        if (3'h2 == state_cache) begin // @[cache.scala 49:26]
          off <= 4'h0; // @[cache.scala 63:25]
        end else begin
          off <= _GEN_515;
        end
      end
    end
    if (reset) begin // @[cache.scala 48:30]
      state_cache <= 3'h0; // @[cache.scala 48:30]
    end else if (3'h0 == state_cache) begin // @[cache.scala 49:26]
      if (_T_1) begin // @[cache.scala 51:34]
        if (hit) begin // @[cache.scala 52:35]
          state_cache <= 3'h1;
        end else begin
          state_cache <= 3'h2;
        end
      end else begin
        state_cache <= 3'h0; // @[cache.scala 54:29]
      end
    end else if (3'h1 == state_cache) begin // @[cache.scala 49:26]
      state_cache <= 3'h0; // @[cache.scala 58:25]
    end else if (3'h2 == state_cache) begin // @[cache.scala 49:26]
      state_cache <= _state_cache_T_2; // @[cache.scala 62:25]
    end else begin
      state_cache <= _GEN_514;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_0[initvar] = _RAND_0[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_1[initvar] = _RAND_3[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_2[initvar] = _RAND_6[31:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_3[initvar] = _RAND_9[31:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_4[initvar] = _RAND_12[31:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_5[initvar] = _RAND_15[31:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_6[initvar] = _RAND_18[31:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_7[initvar] = _RAND_21[31:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_8[initvar] = _RAND_24[31:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_9[initvar] = _RAND_27[31:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_10[initvar] = _RAND_30[31:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_11[initvar] = _RAND_33[31:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_12[initvar] = _RAND_36[31:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_13[initvar] = _RAND_39[31:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_14[initvar] = _RAND_42[31:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_0_15[initvar] = _RAND_45[31:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_0[initvar] = _RAND_48[31:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_1[initvar] = _RAND_51[31:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_2[initvar] = _RAND_54[31:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_3[initvar] = _RAND_57[31:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_4[initvar] = _RAND_60[31:0];
  _RAND_63 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_5[initvar] = _RAND_63[31:0];
  _RAND_66 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_6[initvar] = _RAND_66[31:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_7[initvar] = _RAND_69[31:0];
  _RAND_72 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_8[initvar] = _RAND_72[31:0];
  _RAND_75 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_9[initvar] = _RAND_75[31:0];
  _RAND_78 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_10[initvar] = _RAND_78[31:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_11[initvar] = _RAND_81[31:0];
  _RAND_84 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_12[initvar] = _RAND_84[31:0];
  _RAND_87 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_13[initvar] = _RAND_87[31:0];
  _RAND_90 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_14[initvar] = _RAND_90[31:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_1_15[initvar] = _RAND_93[31:0];
  _RAND_96 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_0[initvar] = _RAND_96[31:0];
  _RAND_99 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_1[initvar] = _RAND_99[31:0];
  _RAND_102 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_2[initvar] = _RAND_102[31:0];
  _RAND_105 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_3[initvar] = _RAND_105[31:0];
  _RAND_108 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_4[initvar] = _RAND_108[31:0];
  _RAND_111 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_5[initvar] = _RAND_111[31:0];
  _RAND_114 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_6[initvar] = _RAND_114[31:0];
  _RAND_117 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_7[initvar] = _RAND_117[31:0];
  _RAND_120 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_8[initvar] = _RAND_120[31:0];
  _RAND_123 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_9[initvar] = _RAND_123[31:0];
  _RAND_126 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_10[initvar] = _RAND_126[31:0];
  _RAND_129 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_11[initvar] = _RAND_129[31:0];
  _RAND_132 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_12[initvar] = _RAND_132[31:0];
  _RAND_135 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_13[initvar] = _RAND_135[31:0];
  _RAND_138 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_14[initvar] = _RAND_138[31:0];
  _RAND_141 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_2_15[initvar] = _RAND_141[31:0];
  _RAND_144 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_0[initvar] = _RAND_144[31:0];
  _RAND_147 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_1[initvar] = _RAND_147[31:0];
  _RAND_150 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_2[initvar] = _RAND_150[31:0];
  _RAND_153 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_3[initvar] = _RAND_153[31:0];
  _RAND_156 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_4[initvar] = _RAND_156[31:0];
  _RAND_159 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_5[initvar] = _RAND_159[31:0];
  _RAND_162 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_6[initvar] = _RAND_162[31:0];
  _RAND_165 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_7[initvar] = _RAND_165[31:0];
  _RAND_168 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_8[initvar] = _RAND_168[31:0];
  _RAND_171 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_9[initvar] = _RAND_171[31:0];
  _RAND_174 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_10[initvar] = _RAND_174[31:0];
  _RAND_177 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_11[initvar] = _RAND_177[31:0];
  _RAND_180 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_12[initvar] = _RAND_180[31:0];
  _RAND_183 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_13[initvar] = _RAND_183[31:0];
  _RAND_186 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_14[initvar] = _RAND_186[31:0];
  _RAND_189 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_3_15[initvar] = _RAND_189[31:0];
  _RAND_192 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_0[initvar] = _RAND_192[31:0];
  _RAND_195 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_1[initvar] = _RAND_195[31:0];
  _RAND_198 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_2[initvar] = _RAND_198[31:0];
  _RAND_201 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_3[initvar] = _RAND_201[31:0];
  _RAND_204 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_4[initvar] = _RAND_204[31:0];
  _RAND_207 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_5[initvar] = _RAND_207[31:0];
  _RAND_210 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_6[initvar] = _RAND_210[31:0];
  _RAND_213 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_7[initvar] = _RAND_213[31:0];
  _RAND_216 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_8[initvar] = _RAND_216[31:0];
  _RAND_219 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_9[initvar] = _RAND_219[31:0];
  _RAND_222 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_10[initvar] = _RAND_222[31:0];
  _RAND_225 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_11[initvar] = _RAND_225[31:0];
  _RAND_228 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_12[initvar] = _RAND_228[31:0];
  _RAND_231 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_13[initvar] = _RAND_231[31:0];
  _RAND_234 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_14[initvar] = _RAND_234[31:0];
  _RAND_237 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_4_15[initvar] = _RAND_237[31:0];
  _RAND_240 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_0[initvar] = _RAND_240[31:0];
  _RAND_243 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_1[initvar] = _RAND_243[31:0];
  _RAND_246 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_2[initvar] = _RAND_246[31:0];
  _RAND_249 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_3[initvar] = _RAND_249[31:0];
  _RAND_252 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_4[initvar] = _RAND_252[31:0];
  _RAND_255 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_5[initvar] = _RAND_255[31:0];
  _RAND_258 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_6[initvar] = _RAND_258[31:0];
  _RAND_261 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_7[initvar] = _RAND_261[31:0];
  _RAND_264 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_8[initvar] = _RAND_264[31:0];
  _RAND_267 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_9[initvar] = _RAND_267[31:0];
  _RAND_270 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_10[initvar] = _RAND_270[31:0];
  _RAND_273 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_11[initvar] = _RAND_273[31:0];
  _RAND_276 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_12[initvar] = _RAND_276[31:0];
  _RAND_279 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_13[initvar] = _RAND_279[31:0];
  _RAND_282 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_14[initvar] = _RAND_282[31:0];
  _RAND_285 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_5_15[initvar] = _RAND_285[31:0];
  _RAND_288 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_0[initvar] = _RAND_288[31:0];
  _RAND_291 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_1[initvar] = _RAND_291[31:0];
  _RAND_294 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_2[initvar] = _RAND_294[31:0];
  _RAND_297 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_3[initvar] = _RAND_297[31:0];
  _RAND_300 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_4[initvar] = _RAND_300[31:0];
  _RAND_303 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_5[initvar] = _RAND_303[31:0];
  _RAND_306 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_6[initvar] = _RAND_306[31:0];
  _RAND_309 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_7[initvar] = _RAND_309[31:0];
  _RAND_312 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_8[initvar] = _RAND_312[31:0];
  _RAND_315 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_9[initvar] = _RAND_315[31:0];
  _RAND_318 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_10[initvar] = _RAND_318[31:0];
  _RAND_321 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_11[initvar] = _RAND_321[31:0];
  _RAND_324 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_12[initvar] = _RAND_324[31:0];
  _RAND_327 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_13[initvar] = _RAND_327[31:0];
  _RAND_330 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_14[initvar] = _RAND_330[31:0];
  _RAND_333 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_6_15[initvar] = _RAND_333[31:0];
  _RAND_336 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_0[initvar] = _RAND_336[31:0];
  _RAND_339 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_1[initvar] = _RAND_339[31:0];
  _RAND_342 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_2[initvar] = _RAND_342[31:0];
  _RAND_345 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_3[initvar] = _RAND_345[31:0];
  _RAND_348 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_4[initvar] = _RAND_348[31:0];
  _RAND_351 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_5[initvar] = _RAND_351[31:0];
  _RAND_354 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_6[initvar] = _RAND_354[31:0];
  _RAND_357 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_7[initvar] = _RAND_357[31:0];
  _RAND_360 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_8[initvar] = _RAND_360[31:0];
  _RAND_363 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_9[initvar] = _RAND_363[31:0];
  _RAND_366 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_10[initvar] = _RAND_366[31:0];
  _RAND_369 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_11[initvar] = _RAND_369[31:0];
  _RAND_372 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_12[initvar] = _RAND_372[31:0];
  _RAND_375 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_13[initvar] = _RAND_375[31:0];
  _RAND_378 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_14[initvar] = _RAND_378[31:0];
  _RAND_381 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_7_15[initvar] = _RAND_381[31:0];
  _RAND_384 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_0[initvar] = _RAND_384[31:0];
  _RAND_387 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_1[initvar] = _RAND_387[31:0];
  _RAND_390 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_2[initvar] = _RAND_390[31:0];
  _RAND_393 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_3[initvar] = _RAND_393[31:0];
  _RAND_396 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_4[initvar] = _RAND_396[31:0];
  _RAND_399 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_5[initvar] = _RAND_399[31:0];
  _RAND_402 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_6[initvar] = _RAND_402[31:0];
  _RAND_405 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_7[initvar] = _RAND_405[31:0];
  _RAND_408 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_8[initvar] = _RAND_408[31:0];
  _RAND_411 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_9[initvar] = _RAND_411[31:0];
  _RAND_414 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_10[initvar] = _RAND_414[31:0];
  _RAND_417 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_11[initvar] = _RAND_417[31:0];
  _RAND_420 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_12[initvar] = _RAND_420[31:0];
  _RAND_423 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_13[initvar] = _RAND_423[31:0];
  _RAND_426 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_14[initvar] = _RAND_426[31:0];
  _RAND_429 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_8_15[initvar] = _RAND_429[31:0];
  _RAND_432 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_0[initvar] = _RAND_432[31:0];
  _RAND_435 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_1[initvar] = _RAND_435[31:0];
  _RAND_438 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_2[initvar] = _RAND_438[31:0];
  _RAND_441 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_3[initvar] = _RAND_441[31:0];
  _RAND_444 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_4[initvar] = _RAND_444[31:0];
  _RAND_447 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_5[initvar] = _RAND_447[31:0];
  _RAND_450 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_6[initvar] = _RAND_450[31:0];
  _RAND_453 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_7[initvar] = _RAND_453[31:0];
  _RAND_456 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_8[initvar] = _RAND_456[31:0];
  _RAND_459 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_9[initvar] = _RAND_459[31:0];
  _RAND_462 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_10[initvar] = _RAND_462[31:0];
  _RAND_465 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_11[initvar] = _RAND_465[31:0];
  _RAND_468 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_12[initvar] = _RAND_468[31:0];
  _RAND_471 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_13[initvar] = _RAND_471[31:0];
  _RAND_474 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_14[initvar] = _RAND_474[31:0];
  _RAND_477 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_9_15[initvar] = _RAND_477[31:0];
  _RAND_480 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_0[initvar] = _RAND_480[31:0];
  _RAND_483 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_1[initvar] = _RAND_483[31:0];
  _RAND_486 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_2[initvar] = _RAND_486[31:0];
  _RAND_489 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_3[initvar] = _RAND_489[31:0];
  _RAND_492 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_4[initvar] = _RAND_492[31:0];
  _RAND_495 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_5[initvar] = _RAND_495[31:0];
  _RAND_498 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_6[initvar] = _RAND_498[31:0];
  _RAND_501 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_7[initvar] = _RAND_501[31:0];
  _RAND_504 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_8[initvar] = _RAND_504[31:0];
  _RAND_507 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_9[initvar] = _RAND_507[31:0];
  _RAND_510 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_10[initvar] = _RAND_510[31:0];
  _RAND_513 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_11[initvar] = _RAND_513[31:0];
  _RAND_516 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_12[initvar] = _RAND_516[31:0];
  _RAND_519 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_13[initvar] = _RAND_519[31:0];
  _RAND_522 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_14[initvar] = _RAND_522[31:0];
  _RAND_525 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_10_15[initvar] = _RAND_525[31:0];
  _RAND_528 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_0[initvar] = _RAND_528[31:0];
  _RAND_531 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_1[initvar] = _RAND_531[31:0];
  _RAND_534 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_2[initvar] = _RAND_534[31:0];
  _RAND_537 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_3[initvar] = _RAND_537[31:0];
  _RAND_540 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_4[initvar] = _RAND_540[31:0];
  _RAND_543 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_5[initvar] = _RAND_543[31:0];
  _RAND_546 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_6[initvar] = _RAND_546[31:0];
  _RAND_549 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_7[initvar] = _RAND_549[31:0];
  _RAND_552 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_8[initvar] = _RAND_552[31:0];
  _RAND_555 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_9[initvar] = _RAND_555[31:0];
  _RAND_558 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_10[initvar] = _RAND_558[31:0];
  _RAND_561 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_11[initvar] = _RAND_561[31:0];
  _RAND_564 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_12[initvar] = _RAND_564[31:0];
  _RAND_567 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_13[initvar] = _RAND_567[31:0];
  _RAND_570 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_14[initvar] = _RAND_570[31:0];
  _RAND_573 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_11_15[initvar] = _RAND_573[31:0];
  _RAND_576 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_0[initvar] = _RAND_576[31:0];
  _RAND_579 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_1[initvar] = _RAND_579[31:0];
  _RAND_582 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_2[initvar] = _RAND_582[31:0];
  _RAND_585 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_3[initvar] = _RAND_585[31:0];
  _RAND_588 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_4[initvar] = _RAND_588[31:0];
  _RAND_591 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_5[initvar] = _RAND_591[31:0];
  _RAND_594 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_6[initvar] = _RAND_594[31:0];
  _RAND_597 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_7[initvar] = _RAND_597[31:0];
  _RAND_600 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_8[initvar] = _RAND_600[31:0];
  _RAND_603 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_9[initvar] = _RAND_603[31:0];
  _RAND_606 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_10[initvar] = _RAND_606[31:0];
  _RAND_609 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_11[initvar] = _RAND_609[31:0];
  _RAND_612 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_12[initvar] = _RAND_612[31:0];
  _RAND_615 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_13[initvar] = _RAND_615[31:0];
  _RAND_618 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_14[initvar] = _RAND_618[31:0];
  _RAND_621 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_12_15[initvar] = _RAND_621[31:0];
  _RAND_624 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_0[initvar] = _RAND_624[31:0];
  _RAND_627 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_1[initvar] = _RAND_627[31:0];
  _RAND_630 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_2[initvar] = _RAND_630[31:0];
  _RAND_633 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_3[initvar] = _RAND_633[31:0];
  _RAND_636 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_4[initvar] = _RAND_636[31:0];
  _RAND_639 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_5[initvar] = _RAND_639[31:0];
  _RAND_642 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_6[initvar] = _RAND_642[31:0];
  _RAND_645 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_7[initvar] = _RAND_645[31:0];
  _RAND_648 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_8[initvar] = _RAND_648[31:0];
  _RAND_651 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_9[initvar] = _RAND_651[31:0];
  _RAND_654 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_10[initvar] = _RAND_654[31:0];
  _RAND_657 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_11[initvar] = _RAND_657[31:0];
  _RAND_660 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_12[initvar] = _RAND_660[31:0];
  _RAND_663 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_13[initvar] = _RAND_663[31:0];
  _RAND_666 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_14[initvar] = _RAND_666[31:0];
  _RAND_669 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_13_15[initvar] = _RAND_669[31:0];
  _RAND_672 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_0[initvar] = _RAND_672[31:0];
  _RAND_675 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_1[initvar] = _RAND_675[31:0];
  _RAND_678 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_2[initvar] = _RAND_678[31:0];
  _RAND_681 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_3[initvar] = _RAND_681[31:0];
  _RAND_684 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_4[initvar] = _RAND_684[31:0];
  _RAND_687 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_5[initvar] = _RAND_687[31:0];
  _RAND_690 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_6[initvar] = _RAND_690[31:0];
  _RAND_693 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_7[initvar] = _RAND_693[31:0];
  _RAND_696 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_8[initvar] = _RAND_696[31:0];
  _RAND_699 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_9[initvar] = _RAND_699[31:0];
  _RAND_702 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_10[initvar] = _RAND_702[31:0];
  _RAND_705 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_11[initvar] = _RAND_705[31:0];
  _RAND_708 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_12[initvar] = _RAND_708[31:0];
  _RAND_711 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_13[initvar] = _RAND_711[31:0];
  _RAND_714 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_14[initvar] = _RAND_714[31:0];
  _RAND_717 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_14_15[initvar] = _RAND_717[31:0];
  _RAND_720 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_0[initvar] = _RAND_720[31:0];
  _RAND_723 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_1[initvar] = _RAND_723[31:0];
  _RAND_726 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_2[initvar] = _RAND_726[31:0];
  _RAND_729 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_3[initvar] = _RAND_729[31:0];
  _RAND_732 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_4[initvar] = _RAND_732[31:0];
  _RAND_735 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_5[initvar] = _RAND_735[31:0];
  _RAND_738 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_6[initvar] = _RAND_738[31:0];
  _RAND_741 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_7[initvar] = _RAND_741[31:0];
  _RAND_744 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_8[initvar] = _RAND_744[31:0];
  _RAND_747 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_9[initvar] = _RAND_747[31:0];
  _RAND_750 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_10[initvar] = _RAND_750[31:0];
  _RAND_753 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_11[initvar] = _RAND_753[31:0];
  _RAND_756 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_12[initvar] = _RAND_756[31:0];
  _RAND_759 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_13[initvar] = _RAND_759[31:0];
  _RAND_762 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_14[initvar] = _RAND_762[31:0];
  _RAND_765 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_15_15[initvar] = _RAND_765[31:0];
  _RAND_768 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_0[initvar] = _RAND_768[31:0];
  _RAND_771 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_1[initvar] = _RAND_771[31:0];
  _RAND_774 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_2[initvar] = _RAND_774[31:0];
  _RAND_777 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_3[initvar] = _RAND_777[31:0];
  _RAND_780 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_4[initvar] = _RAND_780[31:0];
  _RAND_783 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_5[initvar] = _RAND_783[31:0];
  _RAND_786 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_6[initvar] = _RAND_786[31:0];
  _RAND_789 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_7[initvar] = _RAND_789[31:0];
  _RAND_792 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_8[initvar] = _RAND_792[31:0];
  _RAND_795 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_9[initvar] = _RAND_795[31:0];
  _RAND_798 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_10[initvar] = _RAND_798[31:0];
  _RAND_801 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_11[initvar] = _RAND_801[31:0];
  _RAND_804 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_12[initvar] = _RAND_804[31:0];
  _RAND_807 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_13[initvar] = _RAND_807[31:0];
  _RAND_810 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_14[initvar] = _RAND_810[31:0];
  _RAND_813 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_16_15[initvar] = _RAND_813[31:0];
  _RAND_816 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_0[initvar] = _RAND_816[31:0];
  _RAND_819 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_1[initvar] = _RAND_819[31:0];
  _RAND_822 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_2[initvar] = _RAND_822[31:0];
  _RAND_825 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_3[initvar] = _RAND_825[31:0];
  _RAND_828 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_4[initvar] = _RAND_828[31:0];
  _RAND_831 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_5[initvar] = _RAND_831[31:0];
  _RAND_834 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_6[initvar] = _RAND_834[31:0];
  _RAND_837 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_7[initvar] = _RAND_837[31:0];
  _RAND_840 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_8[initvar] = _RAND_840[31:0];
  _RAND_843 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_9[initvar] = _RAND_843[31:0];
  _RAND_846 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_10[initvar] = _RAND_846[31:0];
  _RAND_849 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_11[initvar] = _RAND_849[31:0];
  _RAND_852 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_12[initvar] = _RAND_852[31:0];
  _RAND_855 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_13[initvar] = _RAND_855[31:0];
  _RAND_858 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_14[initvar] = _RAND_858[31:0];
  _RAND_861 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_17_15[initvar] = _RAND_861[31:0];
  _RAND_864 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_0[initvar] = _RAND_864[31:0];
  _RAND_867 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_1[initvar] = _RAND_867[31:0];
  _RAND_870 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_2[initvar] = _RAND_870[31:0];
  _RAND_873 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_3[initvar] = _RAND_873[31:0];
  _RAND_876 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_4[initvar] = _RAND_876[31:0];
  _RAND_879 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_5[initvar] = _RAND_879[31:0];
  _RAND_882 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_6[initvar] = _RAND_882[31:0];
  _RAND_885 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_7[initvar] = _RAND_885[31:0];
  _RAND_888 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_8[initvar] = _RAND_888[31:0];
  _RAND_891 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_9[initvar] = _RAND_891[31:0];
  _RAND_894 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_10[initvar] = _RAND_894[31:0];
  _RAND_897 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_11[initvar] = _RAND_897[31:0];
  _RAND_900 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_12[initvar] = _RAND_900[31:0];
  _RAND_903 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_13[initvar] = _RAND_903[31:0];
  _RAND_906 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_14[initvar] = _RAND_906[31:0];
  _RAND_909 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_18_15[initvar] = _RAND_909[31:0];
  _RAND_912 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_0[initvar] = _RAND_912[31:0];
  _RAND_915 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_1[initvar] = _RAND_915[31:0];
  _RAND_918 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_2[initvar] = _RAND_918[31:0];
  _RAND_921 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_3[initvar] = _RAND_921[31:0];
  _RAND_924 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_4[initvar] = _RAND_924[31:0];
  _RAND_927 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_5[initvar] = _RAND_927[31:0];
  _RAND_930 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_6[initvar] = _RAND_930[31:0];
  _RAND_933 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_7[initvar] = _RAND_933[31:0];
  _RAND_936 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_8[initvar] = _RAND_936[31:0];
  _RAND_939 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_9[initvar] = _RAND_939[31:0];
  _RAND_942 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_10[initvar] = _RAND_942[31:0];
  _RAND_945 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_11[initvar] = _RAND_945[31:0];
  _RAND_948 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_12[initvar] = _RAND_948[31:0];
  _RAND_951 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_13[initvar] = _RAND_951[31:0];
  _RAND_954 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_14[initvar] = _RAND_954[31:0];
  _RAND_957 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_19_15[initvar] = _RAND_957[31:0];
  _RAND_960 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_0[initvar] = _RAND_960[31:0];
  _RAND_963 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_1[initvar] = _RAND_963[31:0];
  _RAND_966 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_2[initvar] = _RAND_966[31:0];
  _RAND_969 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_3[initvar] = _RAND_969[31:0];
  _RAND_972 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_4[initvar] = _RAND_972[31:0];
  _RAND_975 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_5[initvar] = _RAND_975[31:0];
  _RAND_978 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_6[initvar] = _RAND_978[31:0];
  _RAND_981 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_7[initvar] = _RAND_981[31:0];
  _RAND_984 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_8[initvar] = _RAND_984[31:0];
  _RAND_987 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_9[initvar] = _RAND_987[31:0];
  _RAND_990 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_10[initvar] = _RAND_990[31:0];
  _RAND_993 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_11[initvar] = _RAND_993[31:0];
  _RAND_996 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_12[initvar] = _RAND_996[31:0];
  _RAND_999 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_13[initvar] = _RAND_999[31:0];
  _RAND_1002 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_14[initvar] = _RAND_1002[31:0];
  _RAND_1005 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_20_15[initvar] = _RAND_1005[31:0];
  _RAND_1008 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_0[initvar] = _RAND_1008[31:0];
  _RAND_1011 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_1[initvar] = _RAND_1011[31:0];
  _RAND_1014 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_2[initvar] = _RAND_1014[31:0];
  _RAND_1017 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_3[initvar] = _RAND_1017[31:0];
  _RAND_1020 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_4[initvar] = _RAND_1020[31:0];
  _RAND_1023 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_5[initvar] = _RAND_1023[31:0];
  _RAND_1026 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_6[initvar] = _RAND_1026[31:0];
  _RAND_1029 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_7[initvar] = _RAND_1029[31:0];
  _RAND_1032 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_8[initvar] = _RAND_1032[31:0];
  _RAND_1035 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_9[initvar] = _RAND_1035[31:0];
  _RAND_1038 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_10[initvar] = _RAND_1038[31:0];
  _RAND_1041 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_11[initvar] = _RAND_1041[31:0];
  _RAND_1044 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_12[initvar] = _RAND_1044[31:0];
  _RAND_1047 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_13[initvar] = _RAND_1047[31:0];
  _RAND_1050 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_14[initvar] = _RAND_1050[31:0];
  _RAND_1053 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_21_15[initvar] = _RAND_1053[31:0];
  _RAND_1056 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_0[initvar] = _RAND_1056[31:0];
  _RAND_1059 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_1[initvar] = _RAND_1059[31:0];
  _RAND_1062 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_2[initvar] = _RAND_1062[31:0];
  _RAND_1065 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_3[initvar] = _RAND_1065[31:0];
  _RAND_1068 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_4[initvar] = _RAND_1068[31:0];
  _RAND_1071 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_5[initvar] = _RAND_1071[31:0];
  _RAND_1074 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_6[initvar] = _RAND_1074[31:0];
  _RAND_1077 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_7[initvar] = _RAND_1077[31:0];
  _RAND_1080 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_8[initvar] = _RAND_1080[31:0];
  _RAND_1083 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_9[initvar] = _RAND_1083[31:0];
  _RAND_1086 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_10[initvar] = _RAND_1086[31:0];
  _RAND_1089 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_11[initvar] = _RAND_1089[31:0];
  _RAND_1092 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_12[initvar] = _RAND_1092[31:0];
  _RAND_1095 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_13[initvar] = _RAND_1095[31:0];
  _RAND_1098 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_14[initvar] = _RAND_1098[31:0];
  _RAND_1101 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_22_15[initvar] = _RAND_1101[31:0];
  _RAND_1104 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_0[initvar] = _RAND_1104[31:0];
  _RAND_1107 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_1[initvar] = _RAND_1107[31:0];
  _RAND_1110 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_2[initvar] = _RAND_1110[31:0];
  _RAND_1113 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_3[initvar] = _RAND_1113[31:0];
  _RAND_1116 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_4[initvar] = _RAND_1116[31:0];
  _RAND_1119 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_5[initvar] = _RAND_1119[31:0];
  _RAND_1122 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_6[initvar] = _RAND_1122[31:0];
  _RAND_1125 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_7[initvar] = _RAND_1125[31:0];
  _RAND_1128 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_8[initvar] = _RAND_1128[31:0];
  _RAND_1131 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_9[initvar] = _RAND_1131[31:0];
  _RAND_1134 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_10[initvar] = _RAND_1134[31:0];
  _RAND_1137 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_11[initvar] = _RAND_1137[31:0];
  _RAND_1140 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_12[initvar] = _RAND_1140[31:0];
  _RAND_1143 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_13[initvar] = _RAND_1143[31:0];
  _RAND_1146 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_14[initvar] = _RAND_1146[31:0];
  _RAND_1149 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_23_15[initvar] = _RAND_1149[31:0];
  _RAND_1152 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_0[initvar] = _RAND_1152[31:0];
  _RAND_1155 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_1[initvar] = _RAND_1155[31:0];
  _RAND_1158 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_2[initvar] = _RAND_1158[31:0];
  _RAND_1161 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_3[initvar] = _RAND_1161[31:0];
  _RAND_1164 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_4[initvar] = _RAND_1164[31:0];
  _RAND_1167 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_5[initvar] = _RAND_1167[31:0];
  _RAND_1170 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_6[initvar] = _RAND_1170[31:0];
  _RAND_1173 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_7[initvar] = _RAND_1173[31:0];
  _RAND_1176 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_8[initvar] = _RAND_1176[31:0];
  _RAND_1179 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_9[initvar] = _RAND_1179[31:0];
  _RAND_1182 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_10[initvar] = _RAND_1182[31:0];
  _RAND_1185 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_11[initvar] = _RAND_1185[31:0];
  _RAND_1188 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_12[initvar] = _RAND_1188[31:0];
  _RAND_1191 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_13[initvar] = _RAND_1191[31:0];
  _RAND_1194 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_14[initvar] = _RAND_1194[31:0];
  _RAND_1197 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_24_15[initvar] = _RAND_1197[31:0];
  _RAND_1200 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_0[initvar] = _RAND_1200[31:0];
  _RAND_1203 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_1[initvar] = _RAND_1203[31:0];
  _RAND_1206 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_2[initvar] = _RAND_1206[31:0];
  _RAND_1209 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_3[initvar] = _RAND_1209[31:0];
  _RAND_1212 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_4[initvar] = _RAND_1212[31:0];
  _RAND_1215 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_5[initvar] = _RAND_1215[31:0];
  _RAND_1218 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_6[initvar] = _RAND_1218[31:0];
  _RAND_1221 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_7[initvar] = _RAND_1221[31:0];
  _RAND_1224 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_8[initvar] = _RAND_1224[31:0];
  _RAND_1227 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_9[initvar] = _RAND_1227[31:0];
  _RAND_1230 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_10[initvar] = _RAND_1230[31:0];
  _RAND_1233 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_11[initvar] = _RAND_1233[31:0];
  _RAND_1236 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_12[initvar] = _RAND_1236[31:0];
  _RAND_1239 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_13[initvar] = _RAND_1239[31:0];
  _RAND_1242 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_14[initvar] = _RAND_1242[31:0];
  _RAND_1245 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_25_15[initvar] = _RAND_1245[31:0];
  _RAND_1248 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_0[initvar] = _RAND_1248[31:0];
  _RAND_1251 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_1[initvar] = _RAND_1251[31:0];
  _RAND_1254 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_2[initvar] = _RAND_1254[31:0];
  _RAND_1257 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_3[initvar] = _RAND_1257[31:0];
  _RAND_1260 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_4[initvar] = _RAND_1260[31:0];
  _RAND_1263 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_5[initvar] = _RAND_1263[31:0];
  _RAND_1266 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_6[initvar] = _RAND_1266[31:0];
  _RAND_1269 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_7[initvar] = _RAND_1269[31:0];
  _RAND_1272 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_8[initvar] = _RAND_1272[31:0];
  _RAND_1275 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_9[initvar] = _RAND_1275[31:0];
  _RAND_1278 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_10[initvar] = _RAND_1278[31:0];
  _RAND_1281 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_11[initvar] = _RAND_1281[31:0];
  _RAND_1284 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_12[initvar] = _RAND_1284[31:0];
  _RAND_1287 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_13[initvar] = _RAND_1287[31:0];
  _RAND_1290 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_14[initvar] = _RAND_1290[31:0];
  _RAND_1293 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_26_15[initvar] = _RAND_1293[31:0];
  _RAND_1296 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_0[initvar] = _RAND_1296[31:0];
  _RAND_1299 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_1[initvar] = _RAND_1299[31:0];
  _RAND_1302 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_2[initvar] = _RAND_1302[31:0];
  _RAND_1305 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_3[initvar] = _RAND_1305[31:0];
  _RAND_1308 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_4[initvar] = _RAND_1308[31:0];
  _RAND_1311 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_5[initvar] = _RAND_1311[31:0];
  _RAND_1314 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_6[initvar] = _RAND_1314[31:0];
  _RAND_1317 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_7[initvar] = _RAND_1317[31:0];
  _RAND_1320 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_8[initvar] = _RAND_1320[31:0];
  _RAND_1323 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_9[initvar] = _RAND_1323[31:0];
  _RAND_1326 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_10[initvar] = _RAND_1326[31:0];
  _RAND_1329 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_11[initvar] = _RAND_1329[31:0];
  _RAND_1332 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_12[initvar] = _RAND_1332[31:0];
  _RAND_1335 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_13[initvar] = _RAND_1335[31:0];
  _RAND_1338 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_14[initvar] = _RAND_1338[31:0];
  _RAND_1341 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_27_15[initvar] = _RAND_1341[31:0];
  _RAND_1344 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_0[initvar] = _RAND_1344[31:0];
  _RAND_1347 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_1[initvar] = _RAND_1347[31:0];
  _RAND_1350 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_2[initvar] = _RAND_1350[31:0];
  _RAND_1353 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_3[initvar] = _RAND_1353[31:0];
  _RAND_1356 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_4[initvar] = _RAND_1356[31:0];
  _RAND_1359 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_5[initvar] = _RAND_1359[31:0];
  _RAND_1362 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_6[initvar] = _RAND_1362[31:0];
  _RAND_1365 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_7[initvar] = _RAND_1365[31:0];
  _RAND_1368 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_8[initvar] = _RAND_1368[31:0];
  _RAND_1371 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_9[initvar] = _RAND_1371[31:0];
  _RAND_1374 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_10[initvar] = _RAND_1374[31:0];
  _RAND_1377 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_11[initvar] = _RAND_1377[31:0];
  _RAND_1380 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_12[initvar] = _RAND_1380[31:0];
  _RAND_1383 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_13[initvar] = _RAND_1383[31:0];
  _RAND_1386 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_14[initvar] = _RAND_1386[31:0];
  _RAND_1389 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_28_15[initvar] = _RAND_1389[31:0];
  _RAND_1392 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_0[initvar] = _RAND_1392[31:0];
  _RAND_1395 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_1[initvar] = _RAND_1395[31:0];
  _RAND_1398 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_2[initvar] = _RAND_1398[31:0];
  _RAND_1401 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_3[initvar] = _RAND_1401[31:0];
  _RAND_1404 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_4[initvar] = _RAND_1404[31:0];
  _RAND_1407 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_5[initvar] = _RAND_1407[31:0];
  _RAND_1410 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_6[initvar] = _RAND_1410[31:0];
  _RAND_1413 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_7[initvar] = _RAND_1413[31:0];
  _RAND_1416 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_8[initvar] = _RAND_1416[31:0];
  _RAND_1419 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_9[initvar] = _RAND_1419[31:0];
  _RAND_1422 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_10[initvar] = _RAND_1422[31:0];
  _RAND_1425 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_11[initvar] = _RAND_1425[31:0];
  _RAND_1428 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_12[initvar] = _RAND_1428[31:0];
  _RAND_1431 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_13[initvar] = _RAND_1431[31:0];
  _RAND_1434 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_14[initvar] = _RAND_1434[31:0];
  _RAND_1437 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_29_15[initvar] = _RAND_1437[31:0];
  _RAND_1440 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_0[initvar] = _RAND_1440[31:0];
  _RAND_1443 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_1[initvar] = _RAND_1443[31:0];
  _RAND_1446 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_2[initvar] = _RAND_1446[31:0];
  _RAND_1449 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_3[initvar] = _RAND_1449[31:0];
  _RAND_1452 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_4[initvar] = _RAND_1452[31:0];
  _RAND_1455 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_5[initvar] = _RAND_1455[31:0];
  _RAND_1458 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_6[initvar] = _RAND_1458[31:0];
  _RAND_1461 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_7[initvar] = _RAND_1461[31:0];
  _RAND_1464 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_8[initvar] = _RAND_1464[31:0];
  _RAND_1467 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_9[initvar] = _RAND_1467[31:0];
  _RAND_1470 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_10[initvar] = _RAND_1470[31:0];
  _RAND_1473 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_11[initvar] = _RAND_1473[31:0];
  _RAND_1476 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_12[initvar] = _RAND_1476[31:0];
  _RAND_1479 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_13[initvar] = _RAND_1479[31:0];
  _RAND_1482 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_14[initvar] = _RAND_1482[31:0];
  _RAND_1485 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_30_15[initvar] = _RAND_1485[31:0];
  _RAND_1488 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_0[initvar] = _RAND_1488[31:0];
  _RAND_1491 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_1[initvar] = _RAND_1491[31:0];
  _RAND_1494 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_2[initvar] = _RAND_1494[31:0];
  _RAND_1497 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_3[initvar] = _RAND_1497[31:0];
  _RAND_1500 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_4[initvar] = _RAND_1500[31:0];
  _RAND_1503 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_5[initvar] = _RAND_1503[31:0];
  _RAND_1506 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_6[initvar] = _RAND_1506[31:0];
  _RAND_1509 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_7[initvar] = _RAND_1509[31:0];
  _RAND_1512 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_8[initvar] = _RAND_1512[31:0];
  _RAND_1515 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_9[initvar] = _RAND_1515[31:0];
  _RAND_1518 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_10[initvar] = _RAND_1518[31:0];
  _RAND_1521 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_11[initvar] = _RAND_1521[31:0];
  _RAND_1524 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_12[initvar] = _RAND_1524[31:0];
  _RAND_1527 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_13[initvar] = _RAND_1527[31:0];
  _RAND_1530 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_14[initvar] = _RAND_1530[31:0];
  _RAND_1533 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_31_15[initvar] = _RAND_1533[31:0];
  _RAND_1536 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_0[initvar] = _RAND_1536[31:0];
  _RAND_1539 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_1[initvar] = _RAND_1539[31:0];
  _RAND_1542 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_2[initvar] = _RAND_1542[31:0];
  _RAND_1545 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_3[initvar] = _RAND_1545[31:0];
  _RAND_1548 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_4[initvar] = _RAND_1548[31:0];
  _RAND_1551 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_5[initvar] = _RAND_1551[31:0];
  _RAND_1554 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_6[initvar] = _RAND_1554[31:0];
  _RAND_1557 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_7[initvar] = _RAND_1557[31:0];
  _RAND_1560 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_8[initvar] = _RAND_1560[31:0];
  _RAND_1563 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_9[initvar] = _RAND_1563[31:0];
  _RAND_1566 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_10[initvar] = _RAND_1566[31:0];
  _RAND_1569 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_11[initvar] = _RAND_1569[31:0];
  _RAND_1572 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_12[initvar] = _RAND_1572[31:0];
  _RAND_1575 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_13[initvar] = _RAND_1575[31:0];
  _RAND_1578 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_14[initvar] = _RAND_1578[31:0];
  _RAND_1581 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_32_15[initvar] = _RAND_1581[31:0];
  _RAND_1584 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_0[initvar] = _RAND_1584[31:0];
  _RAND_1587 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_1[initvar] = _RAND_1587[31:0];
  _RAND_1590 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_2[initvar] = _RAND_1590[31:0];
  _RAND_1593 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_3[initvar] = _RAND_1593[31:0];
  _RAND_1596 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_4[initvar] = _RAND_1596[31:0];
  _RAND_1599 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_5[initvar] = _RAND_1599[31:0];
  _RAND_1602 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_6[initvar] = _RAND_1602[31:0];
  _RAND_1605 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_7[initvar] = _RAND_1605[31:0];
  _RAND_1608 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_8[initvar] = _RAND_1608[31:0];
  _RAND_1611 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_9[initvar] = _RAND_1611[31:0];
  _RAND_1614 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_10[initvar] = _RAND_1614[31:0];
  _RAND_1617 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_11[initvar] = _RAND_1617[31:0];
  _RAND_1620 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_12[initvar] = _RAND_1620[31:0];
  _RAND_1623 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_13[initvar] = _RAND_1623[31:0];
  _RAND_1626 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_14[initvar] = _RAND_1626[31:0];
  _RAND_1629 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_33_15[initvar] = _RAND_1629[31:0];
  _RAND_1632 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_0[initvar] = _RAND_1632[31:0];
  _RAND_1635 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_1[initvar] = _RAND_1635[31:0];
  _RAND_1638 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_2[initvar] = _RAND_1638[31:0];
  _RAND_1641 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_3[initvar] = _RAND_1641[31:0];
  _RAND_1644 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_4[initvar] = _RAND_1644[31:0];
  _RAND_1647 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_5[initvar] = _RAND_1647[31:0];
  _RAND_1650 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_6[initvar] = _RAND_1650[31:0];
  _RAND_1653 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_7[initvar] = _RAND_1653[31:0];
  _RAND_1656 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_8[initvar] = _RAND_1656[31:0];
  _RAND_1659 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_9[initvar] = _RAND_1659[31:0];
  _RAND_1662 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_10[initvar] = _RAND_1662[31:0];
  _RAND_1665 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_11[initvar] = _RAND_1665[31:0];
  _RAND_1668 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_12[initvar] = _RAND_1668[31:0];
  _RAND_1671 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_13[initvar] = _RAND_1671[31:0];
  _RAND_1674 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_14[initvar] = _RAND_1674[31:0];
  _RAND_1677 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_34_15[initvar] = _RAND_1677[31:0];
  _RAND_1680 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_0[initvar] = _RAND_1680[31:0];
  _RAND_1683 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_1[initvar] = _RAND_1683[31:0];
  _RAND_1686 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_2[initvar] = _RAND_1686[31:0];
  _RAND_1689 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_3[initvar] = _RAND_1689[31:0];
  _RAND_1692 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_4[initvar] = _RAND_1692[31:0];
  _RAND_1695 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_5[initvar] = _RAND_1695[31:0];
  _RAND_1698 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_6[initvar] = _RAND_1698[31:0];
  _RAND_1701 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_7[initvar] = _RAND_1701[31:0];
  _RAND_1704 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_8[initvar] = _RAND_1704[31:0];
  _RAND_1707 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_9[initvar] = _RAND_1707[31:0];
  _RAND_1710 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_10[initvar] = _RAND_1710[31:0];
  _RAND_1713 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_11[initvar] = _RAND_1713[31:0];
  _RAND_1716 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_12[initvar] = _RAND_1716[31:0];
  _RAND_1719 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_13[initvar] = _RAND_1719[31:0];
  _RAND_1722 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_14[initvar] = _RAND_1722[31:0];
  _RAND_1725 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_35_15[initvar] = _RAND_1725[31:0];
  _RAND_1728 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_0[initvar] = _RAND_1728[31:0];
  _RAND_1731 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_1[initvar] = _RAND_1731[31:0];
  _RAND_1734 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_2[initvar] = _RAND_1734[31:0];
  _RAND_1737 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_3[initvar] = _RAND_1737[31:0];
  _RAND_1740 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_4[initvar] = _RAND_1740[31:0];
  _RAND_1743 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_5[initvar] = _RAND_1743[31:0];
  _RAND_1746 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_6[initvar] = _RAND_1746[31:0];
  _RAND_1749 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_7[initvar] = _RAND_1749[31:0];
  _RAND_1752 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_8[initvar] = _RAND_1752[31:0];
  _RAND_1755 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_9[initvar] = _RAND_1755[31:0];
  _RAND_1758 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_10[initvar] = _RAND_1758[31:0];
  _RAND_1761 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_11[initvar] = _RAND_1761[31:0];
  _RAND_1764 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_12[initvar] = _RAND_1764[31:0];
  _RAND_1767 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_13[initvar] = _RAND_1767[31:0];
  _RAND_1770 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_14[initvar] = _RAND_1770[31:0];
  _RAND_1773 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_36_15[initvar] = _RAND_1773[31:0];
  _RAND_1776 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_0[initvar] = _RAND_1776[31:0];
  _RAND_1779 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_1[initvar] = _RAND_1779[31:0];
  _RAND_1782 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_2[initvar] = _RAND_1782[31:0];
  _RAND_1785 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_3[initvar] = _RAND_1785[31:0];
  _RAND_1788 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_4[initvar] = _RAND_1788[31:0];
  _RAND_1791 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_5[initvar] = _RAND_1791[31:0];
  _RAND_1794 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_6[initvar] = _RAND_1794[31:0];
  _RAND_1797 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_7[initvar] = _RAND_1797[31:0];
  _RAND_1800 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_8[initvar] = _RAND_1800[31:0];
  _RAND_1803 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_9[initvar] = _RAND_1803[31:0];
  _RAND_1806 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_10[initvar] = _RAND_1806[31:0];
  _RAND_1809 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_11[initvar] = _RAND_1809[31:0];
  _RAND_1812 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_12[initvar] = _RAND_1812[31:0];
  _RAND_1815 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_13[initvar] = _RAND_1815[31:0];
  _RAND_1818 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_14[initvar] = _RAND_1818[31:0];
  _RAND_1821 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_37_15[initvar] = _RAND_1821[31:0];
  _RAND_1824 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_0[initvar] = _RAND_1824[31:0];
  _RAND_1827 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_1[initvar] = _RAND_1827[31:0];
  _RAND_1830 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_2[initvar] = _RAND_1830[31:0];
  _RAND_1833 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_3[initvar] = _RAND_1833[31:0];
  _RAND_1836 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_4[initvar] = _RAND_1836[31:0];
  _RAND_1839 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_5[initvar] = _RAND_1839[31:0];
  _RAND_1842 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_6[initvar] = _RAND_1842[31:0];
  _RAND_1845 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_7[initvar] = _RAND_1845[31:0];
  _RAND_1848 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_8[initvar] = _RAND_1848[31:0];
  _RAND_1851 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_9[initvar] = _RAND_1851[31:0];
  _RAND_1854 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_10[initvar] = _RAND_1854[31:0];
  _RAND_1857 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_11[initvar] = _RAND_1857[31:0];
  _RAND_1860 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_12[initvar] = _RAND_1860[31:0];
  _RAND_1863 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_13[initvar] = _RAND_1863[31:0];
  _RAND_1866 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_14[initvar] = _RAND_1866[31:0];
  _RAND_1869 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_38_15[initvar] = _RAND_1869[31:0];
  _RAND_1872 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_0[initvar] = _RAND_1872[31:0];
  _RAND_1875 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_1[initvar] = _RAND_1875[31:0];
  _RAND_1878 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_2[initvar] = _RAND_1878[31:0];
  _RAND_1881 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_3[initvar] = _RAND_1881[31:0];
  _RAND_1884 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_4[initvar] = _RAND_1884[31:0];
  _RAND_1887 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_5[initvar] = _RAND_1887[31:0];
  _RAND_1890 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_6[initvar] = _RAND_1890[31:0];
  _RAND_1893 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_7[initvar] = _RAND_1893[31:0];
  _RAND_1896 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_8[initvar] = _RAND_1896[31:0];
  _RAND_1899 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_9[initvar] = _RAND_1899[31:0];
  _RAND_1902 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_10[initvar] = _RAND_1902[31:0];
  _RAND_1905 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_11[initvar] = _RAND_1905[31:0];
  _RAND_1908 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_12[initvar] = _RAND_1908[31:0];
  _RAND_1911 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_13[initvar] = _RAND_1911[31:0];
  _RAND_1914 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_14[initvar] = _RAND_1914[31:0];
  _RAND_1917 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_39_15[initvar] = _RAND_1917[31:0];
  _RAND_1920 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_0[initvar] = _RAND_1920[31:0];
  _RAND_1923 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_1[initvar] = _RAND_1923[31:0];
  _RAND_1926 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_2[initvar] = _RAND_1926[31:0];
  _RAND_1929 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_3[initvar] = _RAND_1929[31:0];
  _RAND_1932 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_4[initvar] = _RAND_1932[31:0];
  _RAND_1935 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_5[initvar] = _RAND_1935[31:0];
  _RAND_1938 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_6[initvar] = _RAND_1938[31:0];
  _RAND_1941 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_7[initvar] = _RAND_1941[31:0];
  _RAND_1944 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_8[initvar] = _RAND_1944[31:0];
  _RAND_1947 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_9[initvar] = _RAND_1947[31:0];
  _RAND_1950 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_10[initvar] = _RAND_1950[31:0];
  _RAND_1953 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_11[initvar] = _RAND_1953[31:0];
  _RAND_1956 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_12[initvar] = _RAND_1956[31:0];
  _RAND_1959 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_13[initvar] = _RAND_1959[31:0];
  _RAND_1962 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_14[initvar] = _RAND_1962[31:0];
  _RAND_1965 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_40_15[initvar] = _RAND_1965[31:0];
  _RAND_1968 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_0[initvar] = _RAND_1968[31:0];
  _RAND_1971 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_1[initvar] = _RAND_1971[31:0];
  _RAND_1974 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_2[initvar] = _RAND_1974[31:0];
  _RAND_1977 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_3[initvar] = _RAND_1977[31:0];
  _RAND_1980 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_4[initvar] = _RAND_1980[31:0];
  _RAND_1983 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_5[initvar] = _RAND_1983[31:0];
  _RAND_1986 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_6[initvar] = _RAND_1986[31:0];
  _RAND_1989 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_7[initvar] = _RAND_1989[31:0];
  _RAND_1992 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_8[initvar] = _RAND_1992[31:0];
  _RAND_1995 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_9[initvar] = _RAND_1995[31:0];
  _RAND_1998 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_10[initvar] = _RAND_1998[31:0];
  _RAND_2001 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_11[initvar] = _RAND_2001[31:0];
  _RAND_2004 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_12[initvar] = _RAND_2004[31:0];
  _RAND_2007 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_13[initvar] = _RAND_2007[31:0];
  _RAND_2010 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_14[initvar] = _RAND_2010[31:0];
  _RAND_2013 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_41_15[initvar] = _RAND_2013[31:0];
  _RAND_2016 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_0[initvar] = _RAND_2016[31:0];
  _RAND_2019 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_1[initvar] = _RAND_2019[31:0];
  _RAND_2022 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_2[initvar] = _RAND_2022[31:0];
  _RAND_2025 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_3[initvar] = _RAND_2025[31:0];
  _RAND_2028 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_4[initvar] = _RAND_2028[31:0];
  _RAND_2031 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_5[initvar] = _RAND_2031[31:0];
  _RAND_2034 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_6[initvar] = _RAND_2034[31:0];
  _RAND_2037 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_7[initvar] = _RAND_2037[31:0];
  _RAND_2040 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_8[initvar] = _RAND_2040[31:0];
  _RAND_2043 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_9[initvar] = _RAND_2043[31:0];
  _RAND_2046 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_10[initvar] = _RAND_2046[31:0];
  _RAND_2049 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_11[initvar] = _RAND_2049[31:0];
  _RAND_2052 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_12[initvar] = _RAND_2052[31:0];
  _RAND_2055 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_13[initvar] = _RAND_2055[31:0];
  _RAND_2058 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_14[initvar] = _RAND_2058[31:0];
  _RAND_2061 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_42_15[initvar] = _RAND_2061[31:0];
  _RAND_2064 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_0[initvar] = _RAND_2064[31:0];
  _RAND_2067 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_1[initvar] = _RAND_2067[31:0];
  _RAND_2070 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_2[initvar] = _RAND_2070[31:0];
  _RAND_2073 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_3[initvar] = _RAND_2073[31:0];
  _RAND_2076 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_4[initvar] = _RAND_2076[31:0];
  _RAND_2079 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_5[initvar] = _RAND_2079[31:0];
  _RAND_2082 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_6[initvar] = _RAND_2082[31:0];
  _RAND_2085 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_7[initvar] = _RAND_2085[31:0];
  _RAND_2088 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_8[initvar] = _RAND_2088[31:0];
  _RAND_2091 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_9[initvar] = _RAND_2091[31:0];
  _RAND_2094 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_10[initvar] = _RAND_2094[31:0];
  _RAND_2097 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_11[initvar] = _RAND_2097[31:0];
  _RAND_2100 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_12[initvar] = _RAND_2100[31:0];
  _RAND_2103 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_13[initvar] = _RAND_2103[31:0];
  _RAND_2106 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_14[initvar] = _RAND_2106[31:0];
  _RAND_2109 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_43_15[initvar] = _RAND_2109[31:0];
  _RAND_2112 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_0[initvar] = _RAND_2112[31:0];
  _RAND_2115 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_1[initvar] = _RAND_2115[31:0];
  _RAND_2118 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_2[initvar] = _RAND_2118[31:0];
  _RAND_2121 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_3[initvar] = _RAND_2121[31:0];
  _RAND_2124 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_4[initvar] = _RAND_2124[31:0];
  _RAND_2127 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_5[initvar] = _RAND_2127[31:0];
  _RAND_2130 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_6[initvar] = _RAND_2130[31:0];
  _RAND_2133 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_7[initvar] = _RAND_2133[31:0];
  _RAND_2136 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_8[initvar] = _RAND_2136[31:0];
  _RAND_2139 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_9[initvar] = _RAND_2139[31:0];
  _RAND_2142 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_10[initvar] = _RAND_2142[31:0];
  _RAND_2145 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_11[initvar] = _RAND_2145[31:0];
  _RAND_2148 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_12[initvar] = _RAND_2148[31:0];
  _RAND_2151 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_13[initvar] = _RAND_2151[31:0];
  _RAND_2154 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_14[initvar] = _RAND_2154[31:0];
  _RAND_2157 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_44_15[initvar] = _RAND_2157[31:0];
  _RAND_2160 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_0[initvar] = _RAND_2160[31:0];
  _RAND_2163 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_1[initvar] = _RAND_2163[31:0];
  _RAND_2166 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_2[initvar] = _RAND_2166[31:0];
  _RAND_2169 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_3[initvar] = _RAND_2169[31:0];
  _RAND_2172 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_4[initvar] = _RAND_2172[31:0];
  _RAND_2175 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_5[initvar] = _RAND_2175[31:0];
  _RAND_2178 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_6[initvar] = _RAND_2178[31:0];
  _RAND_2181 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_7[initvar] = _RAND_2181[31:0];
  _RAND_2184 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_8[initvar] = _RAND_2184[31:0];
  _RAND_2187 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_9[initvar] = _RAND_2187[31:0];
  _RAND_2190 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_10[initvar] = _RAND_2190[31:0];
  _RAND_2193 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_11[initvar] = _RAND_2193[31:0];
  _RAND_2196 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_12[initvar] = _RAND_2196[31:0];
  _RAND_2199 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_13[initvar] = _RAND_2199[31:0];
  _RAND_2202 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_14[initvar] = _RAND_2202[31:0];
  _RAND_2205 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_45_15[initvar] = _RAND_2205[31:0];
  _RAND_2208 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_0[initvar] = _RAND_2208[31:0];
  _RAND_2211 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_1[initvar] = _RAND_2211[31:0];
  _RAND_2214 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_2[initvar] = _RAND_2214[31:0];
  _RAND_2217 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_3[initvar] = _RAND_2217[31:0];
  _RAND_2220 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_4[initvar] = _RAND_2220[31:0];
  _RAND_2223 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_5[initvar] = _RAND_2223[31:0];
  _RAND_2226 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_6[initvar] = _RAND_2226[31:0];
  _RAND_2229 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_7[initvar] = _RAND_2229[31:0];
  _RAND_2232 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_8[initvar] = _RAND_2232[31:0];
  _RAND_2235 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_9[initvar] = _RAND_2235[31:0];
  _RAND_2238 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_10[initvar] = _RAND_2238[31:0];
  _RAND_2241 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_11[initvar] = _RAND_2241[31:0];
  _RAND_2244 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_12[initvar] = _RAND_2244[31:0];
  _RAND_2247 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_13[initvar] = _RAND_2247[31:0];
  _RAND_2250 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_14[initvar] = _RAND_2250[31:0];
  _RAND_2253 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_46_15[initvar] = _RAND_2253[31:0];
  _RAND_2256 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_0[initvar] = _RAND_2256[31:0];
  _RAND_2259 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_1[initvar] = _RAND_2259[31:0];
  _RAND_2262 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_2[initvar] = _RAND_2262[31:0];
  _RAND_2265 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_3[initvar] = _RAND_2265[31:0];
  _RAND_2268 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_4[initvar] = _RAND_2268[31:0];
  _RAND_2271 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_5[initvar] = _RAND_2271[31:0];
  _RAND_2274 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_6[initvar] = _RAND_2274[31:0];
  _RAND_2277 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_7[initvar] = _RAND_2277[31:0];
  _RAND_2280 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_8[initvar] = _RAND_2280[31:0];
  _RAND_2283 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_9[initvar] = _RAND_2283[31:0];
  _RAND_2286 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_10[initvar] = _RAND_2286[31:0];
  _RAND_2289 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_11[initvar] = _RAND_2289[31:0];
  _RAND_2292 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_12[initvar] = _RAND_2292[31:0];
  _RAND_2295 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_13[initvar] = _RAND_2295[31:0];
  _RAND_2298 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_14[initvar] = _RAND_2298[31:0];
  _RAND_2301 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_47_15[initvar] = _RAND_2301[31:0];
  _RAND_2304 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_0[initvar] = _RAND_2304[31:0];
  _RAND_2307 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_1[initvar] = _RAND_2307[31:0];
  _RAND_2310 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_2[initvar] = _RAND_2310[31:0];
  _RAND_2313 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_3[initvar] = _RAND_2313[31:0];
  _RAND_2316 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_4[initvar] = _RAND_2316[31:0];
  _RAND_2319 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_5[initvar] = _RAND_2319[31:0];
  _RAND_2322 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_6[initvar] = _RAND_2322[31:0];
  _RAND_2325 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_7[initvar] = _RAND_2325[31:0];
  _RAND_2328 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_8[initvar] = _RAND_2328[31:0];
  _RAND_2331 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_9[initvar] = _RAND_2331[31:0];
  _RAND_2334 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_10[initvar] = _RAND_2334[31:0];
  _RAND_2337 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_11[initvar] = _RAND_2337[31:0];
  _RAND_2340 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_12[initvar] = _RAND_2340[31:0];
  _RAND_2343 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_13[initvar] = _RAND_2343[31:0];
  _RAND_2346 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_14[initvar] = _RAND_2346[31:0];
  _RAND_2349 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_48_15[initvar] = _RAND_2349[31:0];
  _RAND_2352 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_0[initvar] = _RAND_2352[31:0];
  _RAND_2355 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_1[initvar] = _RAND_2355[31:0];
  _RAND_2358 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_2[initvar] = _RAND_2358[31:0];
  _RAND_2361 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_3[initvar] = _RAND_2361[31:0];
  _RAND_2364 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_4[initvar] = _RAND_2364[31:0];
  _RAND_2367 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_5[initvar] = _RAND_2367[31:0];
  _RAND_2370 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_6[initvar] = _RAND_2370[31:0];
  _RAND_2373 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_7[initvar] = _RAND_2373[31:0];
  _RAND_2376 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_8[initvar] = _RAND_2376[31:0];
  _RAND_2379 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_9[initvar] = _RAND_2379[31:0];
  _RAND_2382 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_10[initvar] = _RAND_2382[31:0];
  _RAND_2385 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_11[initvar] = _RAND_2385[31:0];
  _RAND_2388 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_12[initvar] = _RAND_2388[31:0];
  _RAND_2391 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_13[initvar] = _RAND_2391[31:0];
  _RAND_2394 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_14[initvar] = _RAND_2394[31:0];
  _RAND_2397 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_49_15[initvar] = _RAND_2397[31:0];
  _RAND_2400 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_0[initvar] = _RAND_2400[31:0];
  _RAND_2403 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_1[initvar] = _RAND_2403[31:0];
  _RAND_2406 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_2[initvar] = _RAND_2406[31:0];
  _RAND_2409 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_3[initvar] = _RAND_2409[31:0];
  _RAND_2412 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_4[initvar] = _RAND_2412[31:0];
  _RAND_2415 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_5[initvar] = _RAND_2415[31:0];
  _RAND_2418 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_6[initvar] = _RAND_2418[31:0];
  _RAND_2421 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_7[initvar] = _RAND_2421[31:0];
  _RAND_2424 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_8[initvar] = _RAND_2424[31:0];
  _RAND_2427 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_9[initvar] = _RAND_2427[31:0];
  _RAND_2430 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_10[initvar] = _RAND_2430[31:0];
  _RAND_2433 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_11[initvar] = _RAND_2433[31:0];
  _RAND_2436 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_12[initvar] = _RAND_2436[31:0];
  _RAND_2439 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_13[initvar] = _RAND_2439[31:0];
  _RAND_2442 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_14[initvar] = _RAND_2442[31:0];
  _RAND_2445 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_50_15[initvar] = _RAND_2445[31:0];
  _RAND_2448 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_0[initvar] = _RAND_2448[31:0];
  _RAND_2451 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_1[initvar] = _RAND_2451[31:0];
  _RAND_2454 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_2[initvar] = _RAND_2454[31:0];
  _RAND_2457 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_3[initvar] = _RAND_2457[31:0];
  _RAND_2460 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_4[initvar] = _RAND_2460[31:0];
  _RAND_2463 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_5[initvar] = _RAND_2463[31:0];
  _RAND_2466 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_6[initvar] = _RAND_2466[31:0];
  _RAND_2469 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_7[initvar] = _RAND_2469[31:0];
  _RAND_2472 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_8[initvar] = _RAND_2472[31:0];
  _RAND_2475 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_9[initvar] = _RAND_2475[31:0];
  _RAND_2478 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_10[initvar] = _RAND_2478[31:0];
  _RAND_2481 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_11[initvar] = _RAND_2481[31:0];
  _RAND_2484 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_12[initvar] = _RAND_2484[31:0];
  _RAND_2487 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_13[initvar] = _RAND_2487[31:0];
  _RAND_2490 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_14[initvar] = _RAND_2490[31:0];
  _RAND_2493 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_51_15[initvar] = _RAND_2493[31:0];
  _RAND_2496 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_0[initvar] = _RAND_2496[31:0];
  _RAND_2499 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_1[initvar] = _RAND_2499[31:0];
  _RAND_2502 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_2[initvar] = _RAND_2502[31:0];
  _RAND_2505 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_3[initvar] = _RAND_2505[31:0];
  _RAND_2508 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_4[initvar] = _RAND_2508[31:0];
  _RAND_2511 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_5[initvar] = _RAND_2511[31:0];
  _RAND_2514 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_6[initvar] = _RAND_2514[31:0];
  _RAND_2517 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_7[initvar] = _RAND_2517[31:0];
  _RAND_2520 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_8[initvar] = _RAND_2520[31:0];
  _RAND_2523 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_9[initvar] = _RAND_2523[31:0];
  _RAND_2526 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_10[initvar] = _RAND_2526[31:0];
  _RAND_2529 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_11[initvar] = _RAND_2529[31:0];
  _RAND_2532 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_12[initvar] = _RAND_2532[31:0];
  _RAND_2535 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_13[initvar] = _RAND_2535[31:0];
  _RAND_2538 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_14[initvar] = _RAND_2538[31:0];
  _RAND_2541 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_52_15[initvar] = _RAND_2541[31:0];
  _RAND_2544 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_0[initvar] = _RAND_2544[31:0];
  _RAND_2547 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_1[initvar] = _RAND_2547[31:0];
  _RAND_2550 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_2[initvar] = _RAND_2550[31:0];
  _RAND_2553 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_3[initvar] = _RAND_2553[31:0];
  _RAND_2556 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_4[initvar] = _RAND_2556[31:0];
  _RAND_2559 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_5[initvar] = _RAND_2559[31:0];
  _RAND_2562 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_6[initvar] = _RAND_2562[31:0];
  _RAND_2565 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_7[initvar] = _RAND_2565[31:0];
  _RAND_2568 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_8[initvar] = _RAND_2568[31:0];
  _RAND_2571 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_9[initvar] = _RAND_2571[31:0];
  _RAND_2574 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_10[initvar] = _RAND_2574[31:0];
  _RAND_2577 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_11[initvar] = _RAND_2577[31:0];
  _RAND_2580 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_12[initvar] = _RAND_2580[31:0];
  _RAND_2583 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_13[initvar] = _RAND_2583[31:0];
  _RAND_2586 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_14[initvar] = _RAND_2586[31:0];
  _RAND_2589 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_53_15[initvar] = _RAND_2589[31:0];
  _RAND_2592 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_0[initvar] = _RAND_2592[31:0];
  _RAND_2595 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_1[initvar] = _RAND_2595[31:0];
  _RAND_2598 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_2[initvar] = _RAND_2598[31:0];
  _RAND_2601 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_3[initvar] = _RAND_2601[31:0];
  _RAND_2604 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_4[initvar] = _RAND_2604[31:0];
  _RAND_2607 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_5[initvar] = _RAND_2607[31:0];
  _RAND_2610 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_6[initvar] = _RAND_2610[31:0];
  _RAND_2613 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_7[initvar] = _RAND_2613[31:0];
  _RAND_2616 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_8[initvar] = _RAND_2616[31:0];
  _RAND_2619 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_9[initvar] = _RAND_2619[31:0];
  _RAND_2622 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_10[initvar] = _RAND_2622[31:0];
  _RAND_2625 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_11[initvar] = _RAND_2625[31:0];
  _RAND_2628 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_12[initvar] = _RAND_2628[31:0];
  _RAND_2631 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_13[initvar] = _RAND_2631[31:0];
  _RAND_2634 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_14[initvar] = _RAND_2634[31:0];
  _RAND_2637 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_54_15[initvar] = _RAND_2637[31:0];
  _RAND_2640 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_0[initvar] = _RAND_2640[31:0];
  _RAND_2643 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_1[initvar] = _RAND_2643[31:0];
  _RAND_2646 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_2[initvar] = _RAND_2646[31:0];
  _RAND_2649 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_3[initvar] = _RAND_2649[31:0];
  _RAND_2652 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_4[initvar] = _RAND_2652[31:0];
  _RAND_2655 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_5[initvar] = _RAND_2655[31:0];
  _RAND_2658 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_6[initvar] = _RAND_2658[31:0];
  _RAND_2661 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_7[initvar] = _RAND_2661[31:0];
  _RAND_2664 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_8[initvar] = _RAND_2664[31:0];
  _RAND_2667 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_9[initvar] = _RAND_2667[31:0];
  _RAND_2670 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_10[initvar] = _RAND_2670[31:0];
  _RAND_2673 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_11[initvar] = _RAND_2673[31:0];
  _RAND_2676 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_12[initvar] = _RAND_2676[31:0];
  _RAND_2679 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_13[initvar] = _RAND_2679[31:0];
  _RAND_2682 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_14[initvar] = _RAND_2682[31:0];
  _RAND_2685 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_55_15[initvar] = _RAND_2685[31:0];
  _RAND_2688 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_0[initvar] = _RAND_2688[31:0];
  _RAND_2691 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_1[initvar] = _RAND_2691[31:0];
  _RAND_2694 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_2[initvar] = _RAND_2694[31:0];
  _RAND_2697 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_3[initvar] = _RAND_2697[31:0];
  _RAND_2700 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_4[initvar] = _RAND_2700[31:0];
  _RAND_2703 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_5[initvar] = _RAND_2703[31:0];
  _RAND_2706 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_6[initvar] = _RAND_2706[31:0];
  _RAND_2709 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_7[initvar] = _RAND_2709[31:0];
  _RAND_2712 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_8[initvar] = _RAND_2712[31:0];
  _RAND_2715 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_9[initvar] = _RAND_2715[31:0];
  _RAND_2718 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_10[initvar] = _RAND_2718[31:0];
  _RAND_2721 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_11[initvar] = _RAND_2721[31:0];
  _RAND_2724 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_12[initvar] = _RAND_2724[31:0];
  _RAND_2727 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_13[initvar] = _RAND_2727[31:0];
  _RAND_2730 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_14[initvar] = _RAND_2730[31:0];
  _RAND_2733 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_56_15[initvar] = _RAND_2733[31:0];
  _RAND_2736 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_0[initvar] = _RAND_2736[31:0];
  _RAND_2739 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_1[initvar] = _RAND_2739[31:0];
  _RAND_2742 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_2[initvar] = _RAND_2742[31:0];
  _RAND_2745 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_3[initvar] = _RAND_2745[31:0];
  _RAND_2748 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_4[initvar] = _RAND_2748[31:0];
  _RAND_2751 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_5[initvar] = _RAND_2751[31:0];
  _RAND_2754 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_6[initvar] = _RAND_2754[31:0];
  _RAND_2757 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_7[initvar] = _RAND_2757[31:0];
  _RAND_2760 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_8[initvar] = _RAND_2760[31:0];
  _RAND_2763 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_9[initvar] = _RAND_2763[31:0];
  _RAND_2766 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_10[initvar] = _RAND_2766[31:0];
  _RAND_2769 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_11[initvar] = _RAND_2769[31:0];
  _RAND_2772 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_12[initvar] = _RAND_2772[31:0];
  _RAND_2775 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_13[initvar] = _RAND_2775[31:0];
  _RAND_2778 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_14[initvar] = _RAND_2778[31:0];
  _RAND_2781 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_57_15[initvar] = _RAND_2781[31:0];
  _RAND_2784 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_0[initvar] = _RAND_2784[31:0];
  _RAND_2787 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_1[initvar] = _RAND_2787[31:0];
  _RAND_2790 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_2[initvar] = _RAND_2790[31:0];
  _RAND_2793 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_3[initvar] = _RAND_2793[31:0];
  _RAND_2796 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_4[initvar] = _RAND_2796[31:0];
  _RAND_2799 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_5[initvar] = _RAND_2799[31:0];
  _RAND_2802 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_6[initvar] = _RAND_2802[31:0];
  _RAND_2805 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_7[initvar] = _RAND_2805[31:0];
  _RAND_2808 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_8[initvar] = _RAND_2808[31:0];
  _RAND_2811 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_9[initvar] = _RAND_2811[31:0];
  _RAND_2814 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_10[initvar] = _RAND_2814[31:0];
  _RAND_2817 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_11[initvar] = _RAND_2817[31:0];
  _RAND_2820 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_12[initvar] = _RAND_2820[31:0];
  _RAND_2823 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_13[initvar] = _RAND_2823[31:0];
  _RAND_2826 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_14[initvar] = _RAND_2826[31:0];
  _RAND_2829 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_58_15[initvar] = _RAND_2829[31:0];
  _RAND_2832 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_0[initvar] = _RAND_2832[31:0];
  _RAND_2835 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_1[initvar] = _RAND_2835[31:0];
  _RAND_2838 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_2[initvar] = _RAND_2838[31:0];
  _RAND_2841 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_3[initvar] = _RAND_2841[31:0];
  _RAND_2844 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_4[initvar] = _RAND_2844[31:0];
  _RAND_2847 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_5[initvar] = _RAND_2847[31:0];
  _RAND_2850 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_6[initvar] = _RAND_2850[31:0];
  _RAND_2853 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_7[initvar] = _RAND_2853[31:0];
  _RAND_2856 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_8[initvar] = _RAND_2856[31:0];
  _RAND_2859 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_9[initvar] = _RAND_2859[31:0];
  _RAND_2862 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_10[initvar] = _RAND_2862[31:0];
  _RAND_2865 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_11[initvar] = _RAND_2865[31:0];
  _RAND_2868 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_12[initvar] = _RAND_2868[31:0];
  _RAND_2871 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_13[initvar] = _RAND_2871[31:0];
  _RAND_2874 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_14[initvar] = _RAND_2874[31:0];
  _RAND_2877 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_59_15[initvar] = _RAND_2877[31:0];
  _RAND_2880 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_0[initvar] = _RAND_2880[31:0];
  _RAND_2883 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_1[initvar] = _RAND_2883[31:0];
  _RAND_2886 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_2[initvar] = _RAND_2886[31:0];
  _RAND_2889 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_3[initvar] = _RAND_2889[31:0];
  _RAND_2892 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_4[initvar] = _RAND_2892[31:0];
  _RAND_2895 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_5[initvar] = _RAND_2895[31:0];
  _RAND_2898 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_6[initvar] = _RAND_2898[31:0];
  _RAND_2901 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_7[initvar] = _RAND_2901[31:0];
  _RAND_2904 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_8[initvar] = _RAND_2904[31:0];
  _RAND_2907 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_9[initvar] = _RAND_2907[31:0];
  _RAND_2910 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_10[initvar] = _RAND_2910[31:0];
  _RAND_2913 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_11[initvar] = _RAND_2913[31:0];
  _RAND_2916 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_12[initvar] = _RAND_2916[31:0];
  _RAND_2919 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_13[initvar] = _RAND_2919[31:0];
  _RAND_2922 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_14[initvar] = _RAND_2922[31:0];
  _RAND_2925 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_60_15[initvar] = _RAND_2925[31:0];
  _RAND_2928 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_0[initvar] = _RAND_2928[31:0];
  _RAND_2931 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_1[initvar] = _RAND_2931[31:0];
  _RAND_2934 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_2[initvar] = _RAND_2934[31:0];
  _RAND_2937 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_3[initvar] = _RAND_2937[31:0];
  _RAND_2940 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_4[initvar] = _RAND_2940[31:0];
  _RAND_2943 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_5[initvar] = _RAND_2943[31:0];
  _RAND_2946 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_6[initvar] = _RAND_2946[31:0];
  _RAND_2949 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_7[initvar] = _RAND_2949[31:0];
  _RAND_2952 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_8[initvar] = _RAND_2952[31:0];
  _RAND_2955 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_9[initvar] = _RAND_2955[31:0];
  _RAND_2958 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_10[initvar] = _RAND_2958[31:0];
  _RAND_2961 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_11[initvar] = _RAND_2961[31:0];
  _RAND_2964 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_12[initvar] = _RAND_2964[31:0];
  _RAND_2967 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_13[initvar] = _RAND_2967[31:0];
  _RAND_2970 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_14[initvar] = _RAND_2970[31:0];
  _RAND_2973 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_61_15[initvar] = _RAND_2973[31:0];
  _RAND_2976 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_0[initvar] = _RAND_2976[31:0];
  _RAND_2979 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_1[initvar] = _RAND_2979[31:0];
  _RAND_2982 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_2[initvar] = _RAND_2982[31:0];
  _RAND_2985 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_3[initvar] = _RAND_2985[31:0];
  _RAND_2988 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_4[initvar] = _RAND_2988[31:0];
  _RAND_2991 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_5[initvar] = _RAND_2991[31:0];
  _RAND_2994 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_6[initvar] = _RAND_2994[31:0];
  _RAND_2997 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_7[initvar] = _RAND_2997[31:0];
  _RAND_3000 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_8[initvar] = _RAND_3000[31:0];
  _RAND_3003 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_9[initvar] = _RAND_3003[31:0];
  _RAND_3006 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_10[initvar] = _RAND_3006[31:0];
  _RAND_3009 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_11[initvar] = _RAND_3009[31:0];
  _RAND_3012 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_12[initvar] = _RAND_3012[31:0];
  _RAND_3015 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_13[initvar] = _RAND_3015[31:0];
  _RAND_3018 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_14[initvar] = _RAND_3018[31:0];
  _RAND_3021 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_62_15[initvar] = _RAND_3021[31:0];
  _RAND_3024 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_0[initvar] = _RAND_3024[31:0];
  _RAND_3027 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_1[initvar] = _RAND_3027[31:0];
  _RAND_3030 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_2[initvar] = _RAND_3030[31:0];
  _RAND_3033 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_3[initvar] = _RAND_3033[31:0];
  _RAND_3036 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_4[initvar] = _RAND_3036[31:0];
  _RAND_3039 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_5[initvar] = _RAND_3039[31:0];
  _RAND_3042 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_6[initvar] = _RAND_3042[31:0];
  _RAND_3045 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_7[initvar] = _RAND_3045[31:0];
  _RAND_3048 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_8[initvar] = _RAND_3048[31:0];
  _RAND_3051 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_9[initvar] = _RAND_3051[31:0];
  _RAND_3054 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_10[initvar] = _RAND_3054[31:0];
  _RAND_3057 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_11[initvar] = _RAND_3057[31:0];
  _RAND_3060 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_12[initvar] = _RAND_3060[31:0];
  _RAND_3063 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_13[initvar] = _RAND_3063[31:0];
  _RAND_3066 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_14[initvar] = _RAND_3066[31:0];
  _RAND_3069 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    dataArray_63_15[initvar] = _RAND_3069[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  dataArray_0_0_cachedata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  dataArray_0_0_cachedata_MPORT_addr_pipe_0 = _RAND_2[1:0];
  _RAND_4 = {1{`RANDOM}};
  dataArray_0_1_cachedata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataArray_0_1_cachedata_MPORT_addr_pipe_0 = _RAND_5[1:0];
  _RAND_7 = {1{`RANDOM}};
  dataArray_0_2_cachedata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataArray_0_2_cachedata_MPORT_addr_pipe_0 = _RAND_8[1:0];
  _RAND_10 = {1{`RANDOM}};
  dataArray_0_3_cachedata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataArray_0_3_cachedata_MPORT_addr_pipe_0 = _RAND_11[1:0];
  _RAND_13 = {1{`RANDOM}};
  dataArray_0_4_cachedata_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataArray_0_4_cachedata_MPORT_addr_pipe_0 = _RAND_14[1:0];
  _RAND_16 = {1{`RANDOM}};
  dataArray_0_5_cachedata_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dataArray_0_5_cachedata_MPORT_addr_pipe_0 = _RAND_17[1:0];
  _RAND_19 = {1{`RANDOM}};
  dataArray_0_6_cachedata_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dataArray_0_6_cachedata_MPORT_addr_pipe_0 = _RAND_20[1:0];
  _RAND_22 = {1{`RANDOM}};
  dataArray_0_7_cachedata_MPORT_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  dataArray_0_7_cachedata_MPORT_addr_pipe_0 = _RAND_23[1:0];
  _RAND_25 = {1{`RANDOM}};
  dataArray_0_8_cachedata_MPORT_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  dataArray_0_8_cachedata_MPORT_addr_pipe_0 = _RAND_26[1:0];
  _RAND_28 = {1{`RANDOM}};
  dataArray_0_9_cachedata_MPORT_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dataArray_0_9_cachedata_MPORT_addr_pipe_0 = _RAND_29[1:0];
  _RAND_31 = {1{`RANDOM}};
  dataArray_0_10_cachedata_MPORT_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataArray_0_10_cachedata_MPORT_addr_pipe_0 = _RAND_32[1:0];
  _RAND_34 = {1{`RANDOM}};
  dataArray_0_11_cachedata_MPORT_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataArray_0_11_cachedata_MPORT_addr_pipe_0 = _RAND_35[1:0];
  _RAND_37 = {1{`RANDOM}};
  dataArray_0_12_cachedata_MPORT_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataArray_0_12_cachedata_MPORT_addr_pipe_0 = _RAND_38[1:0];
  _RAND_40 = {1{`RANDOM}};
  dataArray_0_13_cachedata_MPORT_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dataArray_0_13_cachedata_MPORT_addr_pipe_0 = _RAND_41[1:0];
  _RAND_43 = {1{`RANDOM}};
  dataArray_0_14_cachedata_MPORT_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dataArray_0_14_cachedata_MPORT_addr_pipe_0 = _RAND_44[1:0];
  _RAND_46 = {1{`RANDOM}};
  dataArray_0_15_cachedata_MPORT_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dataArray_0_15_cachedata_MPORT_addr_pipe_0 = _RAND_47[1:0];
  _RAND_49 = {1{`RANDOM}};
  dataArray_1_0_cachedata_MPORT_en_pipe_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dataArray_1_0_cachedata_MPORT_addr_pipe_0 = _RAND_50[1:0];
  _RAND_52 = {1{`RANDOM}};
  dataArray_1_1_cachedata_MPORT_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dataArray_1_1_cachedata_MPORT_addr_pipe_0 = _RAND_53[1:0];
  _RAND_55 = {1{`RANDOM}};
  dataArray_1_2_cachedata_MPORT_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dataArray_1_2_cachedata_MPORT_addr_pipe_0 = _RAND_56[1:0];
  _RAND_58 = {1{`RANDOM}};
  dataArray_1_3_cachedata_MPORT_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dataArray_1_3_cachedata_MPORT_addr_pipe_0 = _RAND_59[1:0];
  _RAND_61 = {1{`RANDOM}};
  dataArray_1_4_cachedata_MPORT_en_pipe_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dataArray_1_4_cachedata_MPORT_addr_pipe_0 = _RAND_62[1:0];
  _RAND_64 = {1{`RANDOM}};
  dataArray_1_5_cachedata_MPORT_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dataArray_1_5_cachedata_MPORT_addr_pipe_0 = _RAND_65[1:0];
  _RAND_67 = {1{`RANDOM}};
  dataArray_1_6_cachedata_MPORT_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dataArray_1_6_cachedata_MPORT_addr_pipe_0 = _RAND_68[1:0];
  _RAND_70 = {1{`RANDOM}};
  dataArray_1_7_cachedata_MPORT_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dataArray_1_7_cachedata_MPORT_addr_pipe_0 = _RAND_71[1:0];
  _RAND_73 = {1{`RANDOM}};
  dataArray_1_8_cachedata_MPORT_en_pipe_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dataArray_1_8_cachedata_MPORT_addr_pipe_0 = _RAND_74[1:0];
  _RAND_76 = {1{`RANDOM}};
  dataArray_1_9_cachedata_MPORT_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dataArray_1_9_cachedata_MPORT_addr_pipe_0 = _RAND_77[1:0];
  _RAND_79 = {1{`RANDOM}};
  dataArray_1_10_cachedata_MPORT_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataArray_1_10_cachedata_MPORT_addr_pipe_0 = _RAND_80[1:0];
  _RAND_82 = {1{`RANDOM}};
  dataArray_1_11_cachedata_MPORT_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dataArray_1_11_cachedata_MPORT_addr_pipe_0 = _RAND_83[1:0];
  _RAND_85 = {1{`RANDOM}};
  dataArray_1_12_cachedata_MPORT_en_pipe_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dataArray_1_12_cachedata_MPORT_addr_pipe_0 = _RAND_86[1:0];
  _RAND_88 = {1{`RANDOM}};
  dataArray_1_13_cachedata_MPORT_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dataArray_1_13_cachedata_MPORT_addr_pipe_0 = _RAND_89[1:0];
  _RAND_91 = {1{`RANDOM}};
  dataArray_1_14_cachedata_MPORT_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dataArray_1_14_cachedata_MPORT_addr_pipe_0 = _RAND_92[1:0];
  _RAND_94 = {1{`RANDOM}};
  dataArray_1_15_cachedata_MPORT_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dataArray_1_15_cachedata_MPORT_addr_pipe_0 = _RAND_95[1:0];
  _RAND_97 = {1{`RANDOM}};
  dataArray_2_0_cachedata_MPORT_en_pipe_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dataArray_2_0_cachedata_MPORT_addr_pipe_0 = _RAND_98[1:0];
  _RAND_100 = {1{`RANDOM}};
  dataArray_2_1_cachedata_MPORT_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dataArray_2_1_cachedata_MPORT_addr_pipe_0 = _RAND_101[1:0];
  _RAND_103 = {1{`RANDOM}};
  dataArray_2_2_cachedata_MPORT_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dataArray_2_2_cachedata_MPORT_addr_pipe_0 = _RAND_104[1:0];
  _RAND_106 = {1{`RANDOM}};
  dataArray_2_3_cachedata_MPORT_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dataArray_2_3_cachedata_MPORT_addr_pipe_0 = _RAND_107[1:0];
  _RAND_109 = {1{`RANDOM}};
  dataArray_2_4_cachedata_MPORT_en_pipe_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dataArray_2_4_cachedata_MPORT_addr_pipe_0 = _RAND_110[1:0];
  _RAND_112 = {1{`RANDOM}};
  dataArray_2_5_cachedata_MPORT_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dataArray_2_5_cachedata_MPORT_addr_pipe_0 = _RAND_113[1:0];
  _RAND_115 = {1{`RANDOM}};
  dataArray_2_6_cachedata_MPORT_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dataArray_2_6_cachedata_MPORT_addr_pipe_0 = _RAND_116[1:0];
  _RAND_118 = {1{`RANDOM}};
  dataArray_2_7_cachedata_MPORT_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dataArray_2_7_cachedata_MPORT_addr_pipe_0 = _RAND_119[1:0];
  _RAND_121 = {1{`RANDOM}};
  dataArray_2_8_cachedata_MPORT_en_pipe_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dataArray_2_8_cachedata_MPORT_addr_pipe_0 = _RAND_122[1:0];
  _RAND_124 = {1{`RANDOM}};
  dataArray_2_9_cachedata_MPORT_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dataArray_2_9_cachedata_MPORT_addr_pipe_0 = _RAND_125[1:0];
  _RAND_127 = {1{`RANDOM}};
  dataArray_2_10_cachedata_MPORT_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dataArray_2_10_cachedata_MPORT_addr_pipe_0 = _RAND_128[1:0];
  _RAND_130 = {1{`RANDOM}};
  dataArray_2_11_cachedata_MPORT_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  dataArray_2_11_cachedata_MPORT_addr_pipe_0 = _RAND_131[1:0];
  _RAND_133 = {1{`RANDOM}};
  dataArray_2_12_cachedata_MPORT_en_pipe_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  dataArray_2_12_cachedata_MPORT_addr_pipe_0 = _RAND_134[1:0];
  _RAND_136 = {1{`RANDOM}};
  dataArray_2_13_cachedata_MPORT_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dataArray_2_13_cachedata_MPORT_addr_pipe_0 = _RAND_137[1:0];
  _RAND_139 = {1{`RANDOM}};
  dataArray_2_14_cachedata_MPORT_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dataArray_2_14_cachedata_MPORT_addr_pipe_0 = _RAND_140[1:0];
  _RAND_142 = {1{`RANDOM}};
  dataArray_2_15_cachedata_MPORT_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dataArray_2_15_cachedata_MPORT_addr_pipe_0 = _RAND_143[1:0];
  _RAND_145 = {1{`RANDOM}};
  dataArray_3_0_cachedata_MPORT_en_pipe_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dataArray_3_0_cachedata_MPORT_addr_pipe_0 = _RAND_146[1:0];
  _RAND_148 = {1{`RANDOM}};
  dataArray_3_1_cachedata_MPORT_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dataArray_3_1_cachedata_MPORT_addr_pipe_0 = _RAND_149[1:0];
  _RAND_151 = {1{`RANDOM}};
  dataArray_3_2_cachedata_MPORT_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dataArray_3_2_cachedata_MPORT_addr_pipe_0 = _RAND_152[1:0];
  _RAND_154 = {1{`RANDOM}};
  dataArray_3_3_cachedata_MPORT_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dataArray_3_3_cachedata_MPORT_addr_pipe_0 = _RAND_155[1:0];
  _RAND_157 = {1{`RANDOM}};
  dataArray_3_4_cachedata_MPORT_en_pipe_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dataArray_3_4_cachedata_MPORT_addr_pipe_0 = _RAND_158[1:0];
  _RAND_160 = {1{`RANDOM}};
  dataArray_3_5_cachedata_MPORT_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dataArray_3_5_cachedata_MPORT_addr_pipe_0 = _RAND_161[1:0];
  _RAND_163 = {1{`RANDOM}};
  dataArray_3_6_cachedata_MPORT_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dataArray_3_6_cachedata_MPORT_addr_pipe_0 = _RAND_164[1:0];
  _RAND_166 = {1{`RANDOM}};
  dataArray_3_7_cachedata_MPORT_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dataArray_3_7_cachedata_MPORT_addr_pipe_0 = _RAND_167[1:0];
  _RAND_169 = {1{`RANDOM}};
  dataArray_3_8_cachedata_MPORT_en_pipe_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dataArray_3_8_cachedata_MPORT_addr_pipe_0 = _RAND_170[1:0];
  _RAND_172 = {1{`RANDOM}};
  dataArray_3_9_cachedata_MPORT_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dataArray_3_9_cachedata_MPORT_addr_pipe_0 = _RAND_173[1:0];
  _RAND_175 = {1{`RANDOM}};
  dataArray_3_10_cachedata_MPORT_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dataArray_3_10_cachedata_MPORT_addr_pipe_0 = _RAND_176[1:0];
  _RAND_178 = {1{`RANDOM}};
  dataArray_3_11_cachedata_MPORT_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dataArray_3_11_cachedata_MPORT_addr_pipe_0 = _RAND_179[1:0];
  _RAND_181 = {1{`RANDOM}};
  dataArray_3_12_cachedata_MPORT_en_pipe_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dataArray_3_12_cachedata_MPORT_addr_pipe_0 = _RAND_182[1:0];
  _RAND_184 = {1{`RANDOM}};
  dataArray_3_13_cachedata_MPORT_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dataArray_3_13_cachedata_MPORT_addr_pipe_0 = _RAND_185[1:0];
  _RAND_187 = {1{`RANDOM}};
  dataArray_3_14_cachedata_MPORT_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dataArray_3_14_cachedata_MPORT_addr_pipe_0 = _RAND_188[1:0];
  _RAND_190 = {1{`RANDOM}};
  dataArray_3_15_cachedata_MPORT_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dataArray_3_15_cachedata_MPORT_addr_pipe_0 = _RAND_191[1:0];
  _RAND_193 = {1{`RANDOM}};
  dataArray_4_0_cachedata_MPORT_en_pipe_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dataArray_4_0_cachedata_MPORT_addr_pipe_0 = _RAND_194[1:0];
  _RAND_196 = {1{`RANDOM}};
  dataArray_4_1_cachedata_MPORT_en_pipe_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dataArray_4_1_cachedata_MPORT_addr_pipe_0 = _RAND_197[1:0];
  _RAND_199 = {1{`RANDOM}};
  dataArray_4_2_cachedata_MPORT_en_pipe_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dataArray_4_2_cachedata_MPORT_addr_pipe_0 = _RAND_200[1:0];
  _RAND_202 = {1{`RANDOM}};
  dataArray_4_3_cachedata_MPORT_en_pipe_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dataArray_4_3_cachedata_MPORT_addr_pipe_0 = _RAND_203[1:0];
  _RAND_205 = {1{`RANDOM}};
  dataArray_4_4_cachedata_MPORT_en_pipe_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dataArray_4_4_cachedata_MPORT_addr_pipe_0 = _RAND_206[1:0];
  _RAND_208 = {1{`RANDOM}};
  dataArray_4_5_cachedata_MPORT_en_pipe_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dataArray_4_5_cachedata_MPORT_addr_pipe_0 = _RAND_209[1:0];
  _RAND_211 = {1{`RANDOM}};
  dataArray_4_6_cachedata_MPORT_en_pipe_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dataArray_4_6_cachedata_MPORT_addr_pipe_0 = _RAND_212[1:0];
  _RAND_214 = {1{`RANDOM}};
  dataArray_4_7_cachedata_MPORT_en_pipe_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dataArray_4_7_cachedata_MPORT_addr_pipe_0 = _RAND_215[1:0];
  _RAND_217 = {1{`RANDOM}};
  dataArray_4_8_cachedata_MPORT_en_pipe_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dataArray_4_8_cachedata_MPORT_addr_pipe_0 = _RAND_218[1:0];
  _RAND_220 = {1{`RANDOM}};
  dataArray_4_9_cachedata_MPORT_en_pipe_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dataArray_4_9_cachedata_MPORT_addr_pipe_0 = _RAND_221[1:0];
  _RAND_223 = {1{`RANDOM}};
  dataArray_4_10_cachedata_MPORT_en_pipe_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dataArray_4_10_cachedata_MPORT_addr_pipe_0 = _RAND_224[1:0];
  _RAND_226 = {1{`RANDOM}};
  dataArray_4_11_cachedata_MPORT_en_pipe_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dataArray_4_11_cachedata_MPORT_addr_pipe_0 = _RAND_227[1:0];
  _RAND_229 = {1{`RANDOM}};
  dataArray_4_12_cachedata_MPORT_en_pipe_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dataArray_4_12_cachedata_MPORT_addr_pipe_0 = _RAND_230[1:0];
  _RAND_232 = {1{`RANDOM}};
  dataArray_4_13_cachedata_MPORT_en_pipe_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dataArray_4_13_cachedata_MPORT_addr_pipe_0 = _RAND_233[1:0];
  _RAND_235 = {1{`RANDOM}};
  dataArray_4_14_cachedata_MPORT_en_pipe_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dataArray_4_14_cachedata_MPORT_addr_pipe_0 = _RAND_236[1:0];
  _RAND_238 = {1{`RANDOM}};
  dataArray_4_15_cachedata_MPORT_en_pipe_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dataArray_4_15_cachedata_MPORT_addr_pipe_0 = _RAND_239[1:0];
  _RAND_241 = {1{`RANDOM}};
  dataArray_5_0_cachedata_MPORT_en_pipe_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dataArray_5_0_cachedata_MPORT_addr_pipe_0 = _RAND_242[1:0];
  _RAND_244 = {1{`RANDOM}};
  dataArray_5_1_cachedata_MPORT_en_pipe_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dataArray_5_1_cachedata_MPORT_addr_pipe_0 = _RAND_245[1:0];
  _RAND_247 = {1{`RANDOM}};
  dataArray_5_2_cachedata_MPORT_en_pipe_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dataArray_5_2_cachedata_MPORT_addr_pipe_0 = _RAND_248[1:0];
  _RAND_250 = {1{`RANDOM}};
  dataArray_5_3_cachedata_MPORT_en_pipe_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dataArray_5_3_cachedata_MPORT_addr_pipe_0 = _RAND_251[1:0];
  _RAND_253 = {1{`RANDOM}};
  dataArray_5_4_cachedata_MPORT_en_pipe_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dataArray_5_4_cachedata_MPORT_addr_pipe_0 = _RAND_254[1:0];
  _RAND_256 = {1{`RANDOM}};
  dataArray_5_5_cachedata_MPORT_en_pipe_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  dataArray_5_5_cachedata_MPORT_addr_pipe_0 = _RAND_257[1:0];
  _RAND_259 = {1{`RANDOM}};
  dataArray_5_6_cachedata_MPORT_en_pipe_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dataArray_5_6_cachedata_MPORT_addr_pipe_0 = _RAND_260[1:0];
  _RAND_262 = {1{`RANDOM}};
  dataArray_5_7_cachedata_MPORT_en_pipe_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  dataArray_5_7_cachedata_MPORT_addr_pipe_0 = _RAND_263[1:0];
  _RAND_265 = {1{`RANDOM}};
  dataArray_5_8_cachedata_MPORT_en_pipe_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  dataArray_5_8_cachedata_MPORT_addr_pipe_0 = _RAND_266[1:0];
  _RAND_268 = {1{`RANDOM}};
  dataArray_5_9_cachedata_MPORT_en_pipe_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  dataArray_5_9_cachedata_MPORT_addr_pipe_0 = _RAND_269[1:0];
  _RAND_271 = {1{`RANDOM}};
  dataArray_5_10_cachedata_MPORT_en_pipe_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  dataArray_5_10_cachedata_MPORT_addr_pipe_0 = _RAND_272[1:0];
  _RAND_274 = {1{`RANDOM}};
  dataArray_5_11_cachedata_MPORT_en_pipe_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  dataArray_5_11_cachedata_MPORT_addr_pipe_0 = _RAND_275[1:0];
  _RAND_277 = {1{`RANDOM}};
  dataArray_5_12_cachedata_MPORT_en_pipe_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  dataArray_5_12_cachedata_MPORT_addr_pipe_0 = _RAND_278[1:0];
  _RAND_280 = {1{`RANDOM}};
  dataArray_5_13_cachedata_MPORT_en_pipe_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  dataArray_5_13_cachedata_MPORT_addr_pipe_0 = _RAND_281[1:0];
  _RAND_283 = {1{`RANDOM}};
  dataArray_5_14_cachedata_MPORT_en_pipe_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  dataArray_5_14_cachedata_MPORT_addr_pipe_0 = _RAND_284[1:0];
  _RAND_286 = {1{`RANDOM}};
  dataArray_5_15_cachedata_MPORT_en_pipe_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  dataArray_5_15_cachedata_MPORT_addr_pipe_0 = _RAND_287[1:0];
  _RAND_289 = {1{`RANDOM}};
  dataArray_6_0_cachedata_MPORT_en_pipe_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  dataArray_6_0_cachedata_MPORT_addr_pipe_0 = _RAND_290[1:0];
  _RAND_292 = {1{`RANDOM}};
  dataArray_6_1_cachedata_MPORT_en_pipe_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  dataArray_6_1_cachedata_MPORT_addr_pipe_0 = _RAND_293[1:0];
  _RAND_295 = {1{`RANDOM}};
  dataArray_6_2_cachedata_MPORT_en_pipe_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  dataArray_6_2_cachedata_MPORT_addr_pipe_0 = _RAND_296[1:0];
  _RAND_298 = {1{`RANDOM}};
  dataArray_6_3_cachedata_MPORT_en_pipe_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  dataArray_6_3_cachedata_MPORT_addr_pipe_0 = _RAND_299[1:0];
  _RAND_301 = {1{`RANDOM}};
  dataArray_6_4_cachedata_MPORT_en_pipe_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  dataArray_6_4_cachedata_MPORT_addr_pipe_0 = _RAND_302[1:0];
  _RAND_304 = {1{`RANDOM}};
  dataArray_6_5_cachedata_MPORT_en_pipe_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  dataArray_6_5_cachedata_MPORT_addr_pipe_0 = _RAND_305[1:0];
  _RAND_307 = {1{`RANDOM}};
  dataArray_6_6_cachedata_MPORT_en_pipe_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  dataArray_6_6_cachedata_MPORT_addr_pipe_0 = _RAND_308[1:0];
  _RAND_310 = {1{`RANDOM}};
  dataArray_6_7_cachedata_MPORT_en_pipe_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  dataArray_6_7_cachedata_MPORT_addr_pipe_0 = _RAND_311[1:0];
  _RAND_313 = {1{`RANDOM}};
  dataArray_6_8_cachedata_MPORT_en_pipe_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  dataArray_6_8_cachedata_MPORT_addr_pipe_0 = _RAND_314[1:0];
  _RAND_316 = {1{`RANDOM}};
  dataArray_6_9_cachedata_MPORT_en_pipe_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  dataArray_6_9_cachedata_MPORT_addr_pipe_0 = _RAND_317[1:0];
  _RAND_319 = {1{`RANDOM}};
  dataArray_6_10_cachedata_MPORT_en_pipe_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  dataArray_6_10_cachedata_MPORT_addr_pipe_0 = _RAND_320[1:0];
  _RAND_322 = {1{`RANDOM}};
  dataArray_6_11_cachedata_MPORT_en_pipe_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  dataArray_6_11_cachedata_MPORT_addr_pipe_0 = _RAND_323[1:0];
  _RAND_325 = {1{`RANDOM}};
  dataArray_6_12_cachedata_MPORT_en_pipe_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  dataArray_6_12_cachedata_MPORT_addr_pipe_0 = _RAND_326[1:0];
  _RAND_328 = {1{`RANDOM}};
  dataArray_6_13_cachedata_MPORT_en_pipe_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  dataArray_6_13_cachedata_MPORT_addr_pipe_0 = _RAND_329[1:0];
  _RAND_331 = {1{`RANDOM}};
  dataArray_6_14_cachedata_MPORT_en_pipe_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  dataArray_6_14_cachedata_MPORT_addr_pipe_0 = _RAND_332[1:0];
  _RAND_334 = {1{`RANDOM}};
  dataArray_6_15_cachedata_MPORT_en_pipe_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  dataArray_6_15_cachedata_MPORT_addr_pipe_0 = _RAND_335[1:0];
  _RAND_337 = {1{`RANDOM}};
  dataArray_7_0_cachedata_MPORT_en_pipe_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dataArray_7_0_cachedata_MPORT_addr_pipe_0 = _RAND_338[1:0];
  _RAND_340 = {1{`RANDOM}};
  dataArray_7_1_cachedata_MPORT_en_pipe_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  dataArray_7_1_cachedata_MPORT_addr_pipe_0 = _RAND_341[1:0];
  _RAND_343 = {1{`RANDOM}};
  dataArray_7_2_cachedata_MPORT_en_pipe_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  dataArray_7_2_cachedata_MPORT_addr_pipe_0 = _RAND_344[1:0];
  _RAND_346 = {1{`RANDOM}};
  dataArray_7_3_cachedata_MPORT_en_pipe_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  dataArray_7_3_cachedata_MPORT_addr_pipe_0 = _RAND_347[1:0];
  _RAND_349 = {1{`RANDOM}};
  dataArray_7_4_cachedata_MPORT_en_pipe_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  dataArray_7_4_cachedata_MPORT_addr_pipe_0 = _RAND_350[1:0];
  _RAND_352 = {1{`RANDOM}};
  dataArray_7_5_cachedata_MPORT_en_pipe_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  dataArray_7_5_cachedata_MPORT_addr_pipe_0 = _RAND_353[1:0];
  _RAND_355 = {1{`RANDOM}};
  dataArray_7_6_cachedata_MPORT_en_pipe_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  dataArray_7_6_cachedata_MPORT_addr_pipe_0 = _RAND_356[1:0];
  _RAND_358 = {1{`RANDOM}};
  dataArray_7_7_cachedata_MPORT_en_pipe_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  dataArray_7_7_cachedata_MPORT_addr_pipe_0 = _RAND_359[1:0];
  _RAND_361 = {1{`RANDOM}};
  dataArray_7_8_cachedata_MPORT_en_pipe_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  dataArray_7_8_cachedata_MPORT_addr_pipe_0 = _RAND_362[1:0];
  _RAND_364 = {1{`RANDOM}};
  dataArray_7_9_cachedata_MPORT_en_pipe_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  dataArray_7_9_cachedata_MPORT_addr_pipe_0 = _RAND_365[1:0];
  _RAND_367 = {1{`RANDOM}};
  dataArray_7_10_cachedata_MPORT_en_pipe_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  dataArray_7_10_cachedata_MPORT_addr_pipe_0 = _RAND_368[1:0];
  _RAND_370 = {1{`RANDOM}};
  dataArray_7_11_cachedata_MPORT_en_pipe_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  dataArray_7_11_cachedata_MPORT_addr_pipe_0 = _RAND_371[1:0];
  _RAND_373 = {1{`RANDOM}};
  dataArray_7_12_cachedata_MPORT_en_pipe_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  dataArray_7_12_cachedata_MPORT_addr_pipe_0 = _RAND_374[1:0];
  _RAND_376 = {1{`RANDOM}};
  dataArray_7_13_cachedata_MPORT_en_pipe_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  dataArray_7_13_cachedata_MPORT_addr_pipe_0 = _RAND_377[1:0];
  _RAND_379 = {1{`RANDOM}};
  dataArray_7_14_cachedata_MPORT_en_pipe_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  dataArray_7_14_cachedata_MPORT_addr_pipe_0 = _RAND_380[1:0];
  _RAND_382 = {1{`RANDOM}};
  dataArray_7_15_cachedata_MPORT_en_pipe_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  dataArray_7_15_cachedata_MPORT_addr_pipe_0 = _RAND_383[1:0];
  _RAND_385 = {1{`RANDOM}};
  dataArray_8_0_cachedata_MPORT_en_pipe_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dataArray_8_0_cachedata_MPORT_addr_pipe_0 = _RAND_386[1:0];
  _RAND_388 = {1{`RANDOM}};
  dataArray_8_1_cachedata_MPORT_en_pipe_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dataArray_8_1_cachedata_MPORT_addr_pipe_0 = _RAND_389[1:0];
  _RAND_391 = {1{`RANDOM}};
  dataArray_8_2_cachedata_MPORT_en_pipe_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dataArray_8_2_cachedata_MPORT_addr_pipe_0 = _RAND_392[1:0];
  _RAND_394 = {1{`RANDOM}};
  dataArray_8_3_cachedata_MPORT_en_pipe_0 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dataArray_8_3_cachedata_MPORT_addr_pipe_0 = _RAND_395[1:0];
  _RAND_397 = {1{`RANDOM}};
  dataArray_8_4_cachedata_MPORT_en_pipe_0 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dataArray_8_4_cachedata_MPORT_addr_pipe_0 = _RAND_398[1:0];
  _RAND_400 = {1{`RANDOM}};
  dataArray_8_5_cachedata_MPORT_en_pipe_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dataArray_8_5_cachedata_MPORT_addr_pipe_0 = _RAND_401[1:0];
  _RAND_403 = {1{`RANDOM}};
  dataArray_8_6_cachedata_MPORT_en_pipe_0 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dataArray_8_6_cachedata_MPORT_addr_pipe_0 = _RAND_404[1:0];
  _RAND_406 = {1{`RANDOM}};
  dataArray_8_7_cachedata_MPORT_en_pipe_0 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dataArray_8_7_cachedata_MPORT_addr_pipe_0 = _RAND_407[1:0];
  _RAND_409 = {1{`RANDOM}};
  dataArray_8_8_cachedata_MPORT_en_pipe_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dataArray_8_8_cachedata_MPORT_addr_pipe_0 = _RAND_410[1:0];
  _RAND_412 = {1{`RANDOM}};
  dataArray_8_9_cachedata_MPORT_en_pipe_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dataArray_8_9_cachedata_MPORT_addr_pipe_0 = _RAND_413[1:0];
  _RAND_415 = {1{`RANDOM}};
  dataArray_8_10_cachedata_MPORT_en_pipe_0 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dataArray_8_10_cachedata_MPORT_addr_pipe_0 = _RAND_416[1:0];
  _RAND_418 = {1{`RANDOM}};
  dataArray_8_11_cachedata_MPORT_en_pipe_0 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dataArray_8_11_cachedata_MPORT_addr_pipe_0 = _RAND_419[1:0];
  _RAND_421 = {1{`RANDOM}};
  dataArray_8_12_cachedata_MPORT_en_pipe_0 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dataArray_8_12_cachedata_MPORT_addr_pipe_0 = _RAND_422[1:0];
  _RAND_424 = {1{`RANDOM}};
  dataArray_8_13_cachedata_MPORT_en_pipe_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dataArray_8_13_cachedata_MPORT_addr_pipe_0 = _RAND_425[1:0];
  _RAND_427 = {1{`RANDOM}};
  dataArray_8_14_cachedata_MPORT_en_pipe_0 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dataArray_8_14_cachedata_MPORT_addr_pipe_0 = _RAND_428[1:0];
  _RAND_430 = {1{`RANDOM}};
  dataArray_8_15_cachedata_MPORT_en_pipe_0 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dataArray_8_15_cachedata_MPORT_addr_pipe_0 = _RAND_431[1:0];
  _RAND_433 = {1{`RANDOM}};
  dataArray_9_0_cachedata_MPORT_en_pipe_0 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dataArray_9_0_cachedata_MPORT_addr_pipe_0 = _RAND_434[1:0];
  _RAND_436 = {1{`RANDOM}};
  dataArray_9_1_cachedata_MPORT_en_pipe_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dataArray_9_1_cachedata_MPORT_addr_pipe_0 = _RAND_437[1:0];
  _RAND_439 = {1{`RANDOM}};
  dataArray_9_2_cachedata_MPORT_en_pipe_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dataArray_9_2_cachedata_MPORT_addr_pipe_0 = _RAND_440[1:0];
  _RAND_442 = {1{`RANDOM}};
  dataArray_9_3_cachedata_MPORT_en_pipe_0 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dataArray_9_3_cachedata_MPORT_addr_pipe_0 = _RAND_443[1:0];
  _RAND_445 = {1{`RANDOM}};
  dataArray_9_4_cachedata_MPORT_en_pipe_0 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dataArray_9_4_cachedata_MPORT_addr_pipe_0 = _RAND_446[1:0];
  _RAND_448 = {1{`RANDOM}};
  dataArray_9_5_cachedata_MPORT_en_pipe_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dataArray_9_5_cachedata_MPORT_addr_pipe_0 = _RAND_449[1:0];
  _RAND_451 = {1{`RANDOM}};
  dataArray_9_6_cachedata_MPORT_en_pipe_0 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dataArray_9_6_cachedata_MPORT_addr_pipe_0 = _RAND_452[1:0];
  _RAND_454 = {1{`RANDOM}};
  dataArray_9_7_cachedata_MPORT_en_pipe_0 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dataArray_9_7_cachedata_MPORT_addr_pipe_0 = _RAND_455[1:0];
  _RAND_457 = {1{`RANDOM}};
  dataArray_9_8_cachedata_MPORT_en_pipe_0 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dataArray_9_8_cachedata_MPORT_addr_pipe_0 = _RAND_458[1:0];
  _RAND_460 = {1{`RANDOM}};
  dataArray_9_9_cachedata_MPORT_en_pipe_0 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dataArray_9_9_cachedata_MPORT_addr_pipe_0 = _RAND_461[1:0];
  _RAND_463 = {1{`RANDOM}};
  dataArray_9_10_cachedata_MPORT_en_pipe_0 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dataArray_9_10_cachedata_MPORT_addr_pipe_0 = _RAND_464[1:0];
  _RAND_466 = {1{`RANDOM}};
  dataArray_9_11_cachedata_MPORT_en_pipe_0 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dataArray_9_11_cachedata_MPORT_addr_pipe_0 = _RAND_467[1:0];
  _RAND_469 = {1{`RANDOM}};
  dataArray_9_12_cachedata_MPORT_en_pipe_0 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dataArray_9_12_cachedata_MPORT_addr_pipe_0 = _RAND_470[1:0];
  _RAND_472 = {1{`RANDOM}};
  dataArray_9_13_cachedata_MPORT_en_pipe_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dataArray_9_13_cachedata_MPORT_addr_pipe_0 = _RAND_473[1:0];
  _RAND_475 = {1{`RANDOM}};
  dataArray_9_14_cachedata_MPORT_en_pipe_0 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dataArray_9_14_cachedata_MPORT_addr_pipe_0 = _RAND_476[1:0];
  _RAND_478 = {1{`RANDOM}};
  dataArray_9_15_cachedata_MPORT_en_pipe_0 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dataArray_9_15_cachedata_MPORT_addr_pipe_0 = _RAND_479[1:0];
  _RAND_481 = {1{`RANDOM}};
  dataArray_10_0_cachedata_MPORT_en_pipe_0 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dataArray_10_0_cachedata_MPORT_addr_pipe_0 = _RAND_482[1:0];
  _RAND_484 = {1{`RANDOM}};
  dataArray_10_1_cachedata_MPORT_en_pipe_0 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dataArray_10_1_cachedata_MPORT_addr_pipe_0 = _RAND_485[1:0];
  _RAND_487 = {1{`RANDOM}};
  dataArray_10_2_cachedata_MPORT_en_pipe_0 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dataArray_10_2_cachedata_MPORT_addr_pipe_0 = _RAND_488[1:0];
  _RAND_490 = {1{`RANDOM}};
  dataArray_10_3_cachedata_MPORT_en_pipe_0 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dataArray_10_3_cachedata_MPORT_addr_pipe_0 = _RAND_491[1:0];
  _RAND_493 = {1{`RANDOM}};
  dataArray_10_4_cachedata_MPORT_en_pipe_0 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dataArray_10_4_cachedata_MPORT_addr_pipe_0 = _RAND_494[1:0];
  _RAND_496 = {1{`RANDOM}};
  dataArray_10_5_cachedata_MPORT_en_pipe_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dataArray_10_5_cachedata_MPORT_addr_pipe_0 = _RAND_497[1:0];
  _RAND_499 = {1{`RANDOM}};
  dataArray_10_6_cachedata_MPORT_en_pipe_0 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dataArray_10_6_cachedata_MPORT_addr_pipe_0 = _RAND_500[1:0];
  _RAND_502 = {1{`RANDOM}};
  dataArray_10_7_cachedata_MPORT_en_pipe_0 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dataArray_10_7_cachedata_MPORT_addr_pipe_0 = _RAND_503[1:0];
  _RAND_505 = {1{`RANDOM}};
  dataArray_10_8_cachedata_MPORT_en_pipe_0 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dataArray_10_8_cachedata_MPORT_addr_pipe_0 = _RAND_506[1:0];
  _RAND_508 = {1{`RANDOM}};
  dataArray_10_9_cachedata_MPORT_en_pipe_0 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dataArray_10_9_cachedata_MPORT_addr_pipe_0 = _RAND_509[1:0];
  _RAND_511 = {1{`RANDOM}};
  dataArray_10_10_cachedata_MPORT_en_pipe_0 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dataArray_10_10_cachedata_MPORT_addr_pipe_0 = _RAND_512[1:0];
  _RAND_514 = {1{`RANDOM}};
  dataArray_10_11_cachedata_MPORT_en_pipe_0 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dataArray_10_11_cachedata_MPORT_addr_pipe_0 = _RAND_515[1:0];
  _RAND_517 = {1{`RANDOM}};
  dataArray_10_12_cachedata_MPORT_en_pipe_0 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  dataArray_10_12_cachedata_MPORT_addr_pipe_0 = _RAND_518[1:0];
  _RAND_520 = {1{`RANDOM}};
  dataArray_10_13_cachedata_MPORT_en_pipe_0 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  dataArray_10_13_cachedata_MPORT_addr_pipe_0 = _RAND_521[1:0];
  _RAND_523 = {1{`RANDOM}};
  dataArray_10_14_cachedata_MPORT_en_pipe_0 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  dataArray_10_14_cachedata_MPORT_addr_pipe_0 = _RAND_524[1:0];
  _RAND_526 = {1{`RANDOM}};
  dataArray_10_15_cachedata_MPORT_en_pipe_0 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  dataArray_10_15_cachedata_MPORT_addr_pipe_0 = _RAND_527[1:0];
  _RAND_529 = {1{`RANDOM}};
  dataArray_11_0_cachedata_MPORT_en_pipe_0 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dataArray_11_0_cachedata_MPORT_addr_pipe_0 = _RAND_530[1:0];
  _RAND_532 = {1{`RANDOM}};
  dataArray_11_1_cachedata_MPORT_en_pipe_0 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dataArray_11_1_cachedata_MPORT_addr_pipe_0 = _RAND_533[1:0];
  _RAND_535 = {1{`RANDOM}};
  dataArray_11_2_cachedata_MPORT_en_pipe_0 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  dataArray_11_2_cachedata_MPORT_addr_pipe_0 = _RAND_536[1:0];
  _RAND_538 = {1{`RANDOM}};
  dataArray_11_3_cachedata_MPORT_en_pipe_0 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  dataArray_11_3_cachedata_MPORT_addr_pipe_0 = _RAND_539[1:0];
  _RAND_541 = {1{`RANDOM}};
  dataArray_11_4_cachedata_MPORT_en_pipe_0 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  dataArray_11_4_cachedata_MPORT_addr_pipe_0 = _RAND_542[1:0];
  _RAND_544 = {1{`RANDOM}};
  dataArray_11_5_cachedata_MPORT_en_pipe_0 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  dataArray_11_5_cachedata_MPORT_addr_pipe_0 = _RAND_545[1:0];
  _RAND_547 = {1{`RANDOM}};
  dataArray_11_6_cachedata_MPORT_en_pipe_0 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  dataArray_11_6_cachedata_MPORT_addr_pipe_0 = _RAND_548[1:0];
  _RAND_550 = {1{`RANDOM}};
  dataArray_11_7_cachedata_MPORT_en_pipe_0 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  dataArray_11_7_cachedata_MPORT_addr_pipe_0 = _RAND_551[1:0];
  _RAND_553 = {1{`RANDOM}};
  dataArray_11_8_cachedata_MPORT_en_pipe_0 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dataArray_11_8_cachedata_MPORT_addr_pipe_0 = _RAND_554[1:0];
  _RAND_556 = {1{`RANDOM}};
  dataArray_11_9_cachedata_MPORT_en_pipe_0 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  dataArray_11_9_cachedata_MPORT_addr_pipe_0 = _RAND_557[1:0];
  _RAND_559 = {1{`RANDOM}};
  dataArray_11_10_cachedata_MPORT_en_pipe_0 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  dataArray_11_10_cachedata_MPORT_addr_pipe_0 = _RAND_560[1:0];
  _RAND_562 = {1{`RANDOM}};
  dataArray_11_11_cachedata_MPORT_en_pipe_0 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  dataArray_11_11_cachedata_MPORT_addr_pipe_0 = _RAND_563[1:0];
  _RAND_565 = {1{`RANDOM}};
  dataArray_11_12_cachedata_MPORT_en_pipe_0 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  dataArray_11_12_cachedata_MPORT_addr_pipe_0 = _RAND_566[1:0];
  _RAND_568 = {1{`RANDOM}};
  dataArray_11_13_cachedata_MPORT_en_pipe_0 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  dataArray_11_13_cachedata_MPORT_addr_pipe_0 = _RAND_569[1:0];
  _RAND_571 = {1{`RANDOM}};
  dataArray_11_14_cachedata_MPORT_en_pipe_0 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  dataArray_11_14_cachedata_MPORT_addr_pipe_0 = _RAND_572[1:0];
  _RAND_574 = {1{`RANDOM}};
  dataArray_11_15_cachedata_MPORT_en_pipe_0 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  dataArray_11_15_cachedata_MPORT_addr_pipe_0 = _RAND_575[1:0];
  _RAND_577 = {1{`RANDOM}};
  dataArray_12_0_cachedata_MPORT_en_pipe_0 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  dataArray_12_0_cachedata_MPORT_addr_pipe_0 = _RAND_578[1:0];
  _RAND_580 = {1{`RANDOM}};
  dataArray_12_1_cachedata_MPORT_en_pipe_0 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  dataArray_12_1_cachedata_MPORT_addr_pipe_0 = _RAND_581[1:0];
  _RAND_583 = {1{`RANDOM}};
  dataArray_12_2_cachedata_MPORT_en_pipe_0 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  dataArray_12_2_cachedata_MPORT_addr_pipe_0 = _RAND_584[1:0];
  _RAND_586 = {1{`RANDOM}};
  dataArray_12_3_cachedata_MPORT_en_pipe_0 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  dataArray_12_3_cachedata_MPORT_addr_pipe_0 = _RAND_587[1:0];
  _RAND_589 = {1{`RANDOM}};
  dataArray_12_4_cachedata_MPORT_en_pipe_0 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  dataArray_12_4_cachedata_MPORT_addr_pipe_0 = _RAND_590[1:0];
  _RAND_592 = {1{`RANDOM}};
  dataArray_12_5_cachedata_MPORT_en_pipe_0 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  dataArray_12_5_cachedata_MPORT_addr_pipe_0 = _RAND_593[1:0];
  _RAND_595 = {1{`RANDOM}};
  dataArray_12_6_cachedata_MPORT_en_pipe_0 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  dataArray_12_6_cachedata_MPORT_addr_pipe_0 = _RAND_596[1:0];
  _RAND_598 = {1{`RANDOM}};
  dataArray_12_7_cachedata_MPORT_en_pipe_0 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  dataArray_12_7_cachedata_MPORT_addr_pipe_0 = _RAND_599[1:0];
  _RAND_601 = {1{`RANDOM}};
  dataArray_12_8_cachedata_MPORT_en_pipe_0 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  dataArray_12_8_cachedata_MPORT_addr_pipe_0 = _RAND_602[1:0];
  _RAND_604 = {1{`RANDOM}};
  dataArray_12_9_cachedata_MPORT_en_pipe_0 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  dataArray_12_9_cachedata_MPORT_addr_pipe_0 = _RAND_605[1:0];
  _RAND_607 = {1{`RANDOM}};
  dataArray_12_10_cachedata_MPORT_en_pipe_0 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  dataArray_12_10_cachedata_MPORT_addr_pipe_0 = _RAND_608[1:0];
  _RAND_610 = {1{`RANDOM}};
  dataArray_12_11_cachedata_MPORT_en_pipe_0 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  dataArray_12_11_cachedata_MPORT_addr_pipe_0 = _RAND_611[1:0];
  _RAND_613 = {1{`RANDOM}};
  dataArray_12_12_cachedata_MPORT_en_pipe_0 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  dataArray_12_12_cachedata_MPORT_addr_pipe_0 = _RAND_614[1:0];
  _RAND_616 = {1{`RANDOM}};
  dataArray_12_13_cachedata_MPORT_en_pipe_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  dataArray_12_13_cachedata_MPORT_addr_pipe_0 = _RAND_617[1:0];
  _RAND_619 = {1{`RANDOM}};
  dataArray_12_14_cachedata_MPORT_en_pipe_0 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  dataArray_12_14_cachedata_MPORT_addr_pipe_0 = _RAND_620[1:0];
  _RAND_622 = {1{`RANDOM}};
  dataArray_12_15_cachedata_MPORT_en_pipe_0 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  dataArray_12_15_cachedata_MPORT_addr_pipe_0 = _RAND_623[1:0];
  _RAND_625 = {1{`RANDOM}};
  dataArray_13_0_cachedata_MPORT_en_pipe_0 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  dataArray_13_0_cachedata_MPORT_addr_pipe_0 = _RAND_626[1:0];
  _RAND_628 = {1{`RANDOM}};
  dataArray_13_1_cachedata_MPORT_en_pipe_0 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  dataArray_13_1_cachedata_MPORT_addr_pipe_0 = _RAND_629[1:0];
  _RAND_631 = {1{`RANDOM}};
  dataArray_13_2_cachedata_MPORT_en_pipe_0 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  dataArray_13_2_cachedata_MPORT_addr_pipe_0 = _RAND_632[1:0];
  _RAND_634 = {1{`RANDOM}};
  dataArray_13_3_cachedata_MPORT_en_pipe_0 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  dataArray_13_3_cachedata_MPORT_addr_pipe_0 = _RAND_635[1:0];
  _RAND_637 = {1{`RANDOM}};
  dataArray_13_4_cachedata_MPORT_en_pipe_0 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  dataArray_13_4_cachedata_MPORT_addr_pipe_0 = _RAND_638[1:0];
  _RAND_640 = {1{`RANDOM}};
  dataArray_13_5_cachedata_MPORT_en_pipe_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  dataArray_13_5_cachedata_MPORT_addr_pipe_0 = _RAND_641[1:0];
  _RAND_643 = {1{`RANDOM}};
  dataArray_13_6_cachedata_MPORT_en_pipe_0 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  dataArray_13_6_cachedata_MPORT_addr_pipe_0 = _RAND_644[1:0];
  _RAND_646 = {1{`RANDOM}};
  dataArray_13_7_cachedata_MPORT_en_pipe_0 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  dataArray_13_7_cachedata_MPORT_addr_pipe_0 = _RAND_647[1:0];
  _RAND_649 = {1{`RANDOM}};
  dataArray_13_8_cachedata_MPORT_en_pipe_0 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  dataArray_13_8_cachedata_MPORT_addr_pipe_0 = _RAND_650[1:0];
  _RAND_652 = {1{`RANDOM}};
  dataArray_13_9_cachedata_MPORT_en_pipe_0 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  dataArray_13_9_cachedata_MPORT_addr_pipe_0 = _RAND_653[1:0];
  _RAND_655 = {1{`RANDOM}};
  dataArray_13_10_cachedata_MPORT_en_pipe_0 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  dataArray_13_10_cachedata_MPORT_addr_pipe_0 = _RAND_656[1:0];
  _RAND_658 = {1{`RANDOM}};
  dataArray_13_11_cachedata_MPORT_en_pipe_0 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  dataArray_13_11_cachedata_MPORT_addr_pipe_0 = _RAND_659[1:0];
  _RAND_661 = {1{`RANDOM}};
  dataArray_13_12_cachedata_MPORT_en_pipe_0 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  dataArray_13_12_cachedata_MPORT_addr_pipe_0 = _RAND_662[1:0];
  _RAND_664 = {1{`RANDOM}};
  dataArray_13_13_cachedata_MPORT_en_pipe_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  dataArray_13_13_cachedata_MPORT_addr_pipe_0 = _RAND_665[1:0];
  _RAND_667 = {1{`RANDOM}};
  dataArray_13_14_cachedata_MPORT_en_pipe_0 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  dataArray_13_14_cachedata_MPORT_addr_pipe_0 = _RAND_668[1:0];
  _RAND_670 = {1{`RANDOM}};
  dataArray_13_15_cachedata_MPORT_en_pipe_0 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  dataArray_13_15_cachedata_MPORT_addr_pipe_0 = _RAND_671[1:0];
  _RAND_673 = {1{`RANDOM}};
  dataArray_14_0_cachedata_MPORT_en_pipe_0 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  dataArray_14_0_cachedata_MPORT_addr_pipe_0 = _RAND_674[1:0];
  _RAND_676 = {1{`RANDOM}};
  dataArray_14_1_cachedata_MPORT_en_pipe_0 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  dataArray_14_1_cachedata_MPORT_addr_pipe_0 = _RAND_677[1:0];
  _RAND_679 = {1{`RANDOM}};
  dataArray_14_2_cachedata_MPORT_en_pipe_0 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  dataArray_14_2_cachedata_MPORT_addr_pipe_0 = _RAND_680[1:0];
  _RAND_682 = {1{`RANDOM}};
  dataArray_14_3_cachedata_MPORT_en_pipe_0 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  dataArray_14_3_cachedata_MPORT_addr_pipe_0 = _RAND_683[1:0];
  _RAND_685 = {1{`RANDOM}};
  dataArray_14_4_cachedata_MPORT_en_pipe_0 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  dataArray_14_4_cachedata_MPORT_addr_pipe_0 = _RAND_686[1:0];
  _RAND_688 = {1{`RANDOM}};
  dataArray_14_5_cachedata_MPORT_en_pipe_0 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  dataArray_14_5_cachedata_MPORT_addr_pipe_0 = _RAND_689[1:0];
  _RAND_691 = {1{`RANDOM}};
  dataArray_14_6_cachedata_MPORT_en_pipe_0 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  dataArray_14_6_cachedata_MPORT_addr_pipe_0 = _RAND_692[1:0];
  _RAND_694 = {1{`RANDOM}};
  dataArray_14_7_cachedata_MPORT_en_pipe_0 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  dataArray_14_7_cachedata_MPORT_addr_pipe_0 = _RAND_695[1:0];
  _RAND_697 = {1{`RANDOM}};
  dataArray_14_8_cachedata_MPORT_en_pipe_0 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  dataArray_14_8_cachedata_MPORT_addr_pipe_0 = _RAND_698[1:0];
  _RAND_700 = {1{`RANDOM}};
  dataArray_14_9_cachedata_MPORT_en_pipe_0 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  dataArray_14_9_cachedata_MPORT_addr_pipe_0 = _RAND_701[1:0];
  _RAND_703 = {1{`RANDOM}};
  dataArray_14_10_cachedata_MPORT_en_pipe_0 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  dataArray_14_10_cachedata_MPORT_addr_pipe_0 = _RAND_704[1:0];
  _RAND_706 = {1{`RANDOM}};
  dataArray_14_11_cachedata_MPORT_en_pipe_0 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  dataArray_14_11_cachedata_MPORT_addr_pipe_0 = _RAND_707[1:0];
  _RAND_709 = {1{`RANDOM}};
  dataArray_14_12_cachedata_MPORT_en_pipe_0 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  dataArray_14_12_cachedata_MPORT_addr_pipe_0 = _RAND_710[1:0];
  _RAND_712 = {1{`RANDOM}};
  dataArray_14_13_cachedata_MPORT_en_pipe_0 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  dataArray_14_13_cachedata_MPORT_addr_pipe_0 = _RAND_713[1:0];
  _RAND_715 = {1{`RANDOM}};
  dataArray_14_14_cachedata_MPORT_en_pipe_0 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  dataArray_14_14_cachedata_MPORT_addr_pipe_0 = _RAND_716[1:0];
  _RAND_718 = {1{`RANDOM}};
  dataArray_14_15_cachedata_MPORT_en_pipe_0 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  dataArray_14_15_cachedata_MPORT_addr_pipe_0 = _RAND_719[1:0];
  _RAND_721 = {1{`RANDOM}};
  dataArray_15_0_cachedata_MPORT_en_pipe_0 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  dataArray_15_0_cachedata_MPORT_addr_pipe_0 = _RAND_722[1:0];
  _RAND_724 = {1{`RANDOM}};
  dataArray_15_1_cachedata_MPORT_en_pipe_0 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  dataArray_15_1_cachedata_MPORT_addr_pipe_0 = _RAND_725[1:0];
  _RAND_727 = {1{`RANDOM}};
  dataArray_15_2_cachedata_MPORT_en_pipe_0 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  dataArray_15_2_cachedata_MPORT_addr_pipe_0 = _RAND_728[1:0];
  _RAND_730 = {1{`RANDOM}};
  dataArray_15_3_cachedata_MPORT_en_pipe_0 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  dataArray_15_3_cachedata_MPORT_addr_pipe_0 = _RAND_731[1:0];
  _RAND_733 = {1{`RANDOM}};
  dataArray_15_4_cachedata_MPORT_en_pipe_0 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  dataArray_15_4_cachedata_MPORT_addr_pipe_0 = _RAND_734[1:0];
  _RAND_736 = {1{`RANDOM}};
  dataArray_15_5_cachedata_MPORT_en_pipe_0 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  dataArray_15_5_cachedata_MPORT_addr_pipe_0 = _RAND_737[1:0];
  _RAND_739 = {1{`RANDOM}};
  dataArray_15_6_cachedata_MPORT_en_pipe_0 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  dataArray_15_6_cachedata_MPORT_addr_pipe_0 = _RAND_740[1:0];
  _RAND_742 = {1{`RANDOM}};
  dataArray_15_7_cachedata_MPORT_en_pipe_0 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  dataArray_15_7_cachedata_MPORT_addr_pipe_0 = _RAND_743[1:0];
  _RAND_745 = {1{`RANDOM}};
  dataArray_15_8_cachedata_MPORT_en_pipe_0 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  dataArray_15_8_cachedata_MPORT_addr_pipe_0 = _RAND_746[1:0];
  _RAND_748 = {1{`RANDOM}};
  dataArray_15_9_cachedata_MPORT_en_pipe_0 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  dataArray_15_9_cachedata_MPORT_addr_pipe_0 = _RAND_749[1:0];
  _RAND_751 = {1{`RANDOM}};
  dataArray_15_10_cachedata_MPORT_en_pipe_0 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  dataArray_15_10_cachedata_MPORT_addr_pipe_0 = _RAND_752[1:0];
  _RAND_754 = {1{`RANDOM}};
  dataArray_15_11_cachedata_MPORT_en_pipe_0 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  dataArray_15_11_cachedata_MPORT_addr_pipe_0 = _RAND_755[1:0];
  _RAND_757 = {1{`RANDOM}};
  dataArray_15_12_cachedata_MPORT_en_pipe_0 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  dataArray_15_12_cachedata_MPORT_addr_pipe_0 = _RAND_758[1:0];
  _RAND_760 = {1{`RANDOM}};
  dataArray_15_13_cachedata_MPORT_en_pipe_0 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  dataArray_15_13_cachedata_MPORT_addr_pipe_0 = _RAND_761[1:0];
  _RAND_763 = {1{`RANDOM}};
  dataArray_15_14_cachedata_MPORT_en_pipe_0 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  dataArray_15_14_cachedata_MPORT_addr_pipe_0 = _RAND_764[1:0];
  _RAND_766 = {1{`RANDOM}};
  dataArray_15_15_cachedata_MPORT_en_pipe_0 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  dataArray_15_15_cachedata_MPORT_addr_pipe_0 = _RAND_767[1:0];
  _RAND_769 = {1{`RANDOM}};
  dataArray_16_0_cachedata_MPORT_en_pipe_0 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  dataArray_16_0_cachedata_MPORT_addr_pipe_0 = _RAND_770[1:0];
  _RAND_772 = {1{`RANDOM}};
  dataArray_16_1_cachedata_MPORT_en_pipe_0 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  dataArray_16_1_cachedata_MPORT_addr_pipe_0 = _RAND_773[1:0];
  _RAND_775 = {1{`RANDOM}};
  dataArray_16_2_cachedata_MPORT_en_pipe_0 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  dataArray_16_2_cachedata_MPORT_addr_pipe_0 = _RAND_776[1:0];
  _RAND_778 = {1{`RANDOM}};
  dataArray_16_3_cachedata_MPORT_en_pipe_0 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  dataArray_16_3_cachedata_MPORT_addr_pipe_0 = _RAND_779[1:0];
  _RAND_781 = {1{`RANDOM}};
  dataArray_16_4_cachedata_MPORT_en_pipe_0 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  dataArray_16_4_cachedata_MPORT_addr_pipe_0 = _RAND_782[1:0];
  _RAND_784 = {1{`RANDOM}};
  dataArray_16_5_cachedata_MPORT_en_pipe_0 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  dataArray_16_5_cachedata_MPORT_addr_pipe_0 = _RAND_785[1:0];
  _RAND_787 = {1{`RANDOM}};
  dataArray_16_6_cachedata_MPORT_en_pipe_0 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  dataArray_16_6_cachedata_MPORT_addr_pipe_0 = _RAND_788[1:0];
  _RAND_790 = {1{`RANDOM}};
  dataArray_16_7_cachedata_MPORT_en_pipe_0 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  dataArray_16_7_cachedata_MPORT_addr_pipe_0 = _RAND_791[1:0];
  _RAND_793 = {1{`RANDOM}};
  dataArray_16_8_cachedata_MPORT_en_pipe_0 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  dataArray_16_8_cachedata_MPORT_addr_pipe_0 = _RAND_794[1:0];
  _RAND_796 = {1{`RANDOM}};
  dataArray_16_9_cachedata_MPORT_en_pipe_0 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  dataArray_16_9_cachedata_MPORT_addr_pipe_0 = _RAND_797[1:0];
  _RAND_799 = {1{`RANDOM}};
  dataArray_16_10_cachedata_MPORT_en_pipe_0 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  dataArray_16_10_cachedata_MPORT_addr_pipe_0 = _RAND_800[1:0];
  _RAND_802 = {1{`RANDOM}};
  dataArray_16_11_cachedata_MPORT_en_pipe_0 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  dataArray_16_11_cachedata_MPORT_addr_pipe_0 = _RAND_803[1:0];
  _RAND_805 = {1{`RANDOM}};
  dataArray_16_12_cachedata_MPORT_en_pipe_0 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  dataArray_16_12_cachedata_MPORT_addr_pipe_0 = _RAND_806[1:0];
  _RAND_808 = {1{`RANDOM}};
  dataArray_16_13_cachedata_MPORT_en_pipe_0 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  dataArray_16_13_cachedata_MPORT_addr_pipe_0 = _RAND_809[1:0];
  _RAND_811 = {1{`RANDOM}};
  dataArray_16_14_cachedata_MPORT_en_pipe_0 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  dataArray_16_14_cachedata_MPORT_addr_pipe_0 = _RAND_812[1:0];
  _RAND_814 = {1{`RANDOM}};
  dataArray_16_15_cachedata_MPORT_en_pipe_0 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  dataArray_16_15_cachedata_MPORT_addr_pipe_0 = _RAND_815[1:0];
  _RAND_817 = {1{`RANDOM}};
  dataArray_17_0_cachedata_MPORT_en_pipe_0 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  dataArray_17_0_cachedata_MPORT_addr_pipe_0 = _RAND_818[1:0];
  _RAND_820 = {1{`RANDOM}};
  dataArray_17_1_cachedata_MPORT_en_pipe_0 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  dataArray_17_1_cachedata_MPORT_addr_pipe_0 = _RAND_821[1:0];
  _RAND_823 = {1{`RANDOM}};
  dataArray_17_2_cachedata_MPORT_en_pipe_0 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  dataArray_17_2_cachedata_MPORT_addr_pipe_0 = _RAND_824[1:0];
  _RAND_826 = {1{`RANDOM}};
  dataArray_17_3_cachedata_MPORT_en_pipe_0 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  dataArray_17_3_cachedata_MPORT_addr_pipe_0 = _RAND_827[1:0];
  _RAND_829 = {1{`RANDOM}};
  dataArray_17_4_cachedata_MPORT_en_pipe_0 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  dataArray_17_4_cachedata_MPORT_addr_pipe_0 = _RAND_830[1:0];
  _RAND_832 = {1{`RANDOM}};
  dataArray_17_5_cachedata_MPORT_en_pipe_0 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  dataArray_17_5_cachedata_MPORT_addr_pipe_0 = _RAND_833[1:0];
  _RAND_835 = {1{`RANDOM}};
  dataArray_17_6_cachedata_MPORT_en_pipe_0 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  dataArray_17_6_cachedata_MPORT_addr_pipe_0 = _RAND_836[1:0];
  _RAND_838 = {1{`RANDOM}};
  dataArray_17_7_cachedata_MPORT_en_pipe_0 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  dataArray_17_7_cachedata_MPORT_addr_pipe_0 = _RAND_839[1:0];
  _RAND_841 = {1{`RANDOM}};
  dataArray_17_8_cachedata_MPORT_en_pipe_0 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  dataArray_17_8_cachedata_MPORT_addr_pipe_0 = _RAND_842[1:0];
  _RAND_844 = {1{`RANDOM}};
  dataArray_17_9_cachedata_MPORT_en_pipe_0 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  dataArray_17_9_cachedata_MPORT_addr_pipe_0 = _RAND_845[1:0];
  _RAND_847 = {1{`RANDOM}};
  dataArray_17_10_cachedata_MPORT_en_pipe_0 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  dataArray_17_10_cachedata_MPORT_addr_pipe_0 = _RAND_848[1:0];
  _RAND_850 = {1{`RANDOM}};
  dataArray_17_11_cachedata_MPORT_en_pipe_0 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  dataArray_17_11_cachedata_MPORT_addr_pipe_0 = _RAND_851[1:0];
  _RAND_853 = {1{`RANDOM}};
  dataArray_17_12_cachedata_MPORT_en_pipe_0 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  dataArray_17_12_cachedata_MPORT_addr_pipe_0 = _RAND_854[1:0];
  _RAND_856 = {1{`RANDOM}};
  dataArray_17_13_cachedata_MPORT_en_pipe_0 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  dataArray_17_13_cachedata_MPORT_addr_pipe_0 = _RAND_857[1:0];
  _RAND_859 = {1{`RANDOM}};
  dataArray_17_14_cachedata_MPORT_en_pipe_0 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  dataArray_17_14_cachedata_MPORT_addr_pipe_0 = _RAND_860[1:0];
  _RAND_862 = {1{`RANDOM}};
  dataArray_17_15_cachedata_MPORT_en_pipe_0 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  dataArray_17_15_cachedata_MPORT_addr_pipe_0 = _RAND_863[1:0];
  _RAND_865 = {1{`RANDOM}};
  dataArray_18_0_cachedata_MPORT_en_pipe_0 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  dataArray_18_0_cachedata_MPORT_addr_pipe_0 = _RAND_866[1:0];
  _RAND_868 = {1{`RANDOM}};
  dataArray_18_1_cachedata_MPORT_en_pipe_0 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  dataArray_18_1_cachedata_MPORT_addr_pipe_0 = _RAND_869[1:0];
  _RAND_871 = {1{`RANDOM}};
  dataArray_18_2_cachedata_MPORT_en_pipe_0 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  dataArray_18_2_cachedata_MPORT_addr_pipe_0 = _RAND_872[1:0];
  _RAND_874 = {1{`RANDOM}};
  dataArray_18_3_cachedata_MPORT_en_pipe_0 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  dataArray_18_3_cachedata_MPORT_addr_pipe_0 = _RAND_875[1:0];
  _RAND_877 = {1{`RANDOM}};
  dataArray_18_4_cachedata_MPORT_en_pipe_0 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  dataArray_18_4_cachedata_MPORT_addr_pipe_0 = _RAND_878[1:0];
  _RAND_880 = {1{`RANDOM}};
  dataArray_18_5_cachedata_MPORT_en_pipe_0 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  dataArray_18_5_cachedata_MPORT_addr_pipe_0 = _RAND_881[1:0];
  _RAND_883 = {1{`RANDOM}};
  dataArray_18_6_cachedata_MPORT_en_pipe_0 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  dataArray_18_6_cachedata_MPORT_addr_pipe_0 = _RAND_884[1:0];
  _RAND_886 = {1{`RANDOM}};
  dataArray_18_7_cachedata_MPORT_en_pipe_0 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  dataArray_18_7_cachedata_MPORT_addr_pipe_0 = _RAND_887[1:0];
  _RAND_889 = {1{`RANDOM}};
  dataArray_18_8_cachedata_MPORT_en_pipe_0 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  dataArray_18_8_cachedata_MPORT_addr_pipe_0 = _RAND_890[1:0];
  _RAND_892 = {1{`RANDOM}};
  dataArray_18_9_cachedata_MPORT_en_pipe_0 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  dataArray_18_9_cachedata_MPORT_addr_pipe_0 = _RAND_893[1:0];
  _RAND_895 = {1{`RANDOM}};
  dataArray_18_10_cachedata_MPORT_en_pipe_0 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  dataArray_18_10_cachedata_MPORT_addr_pipe_0 = _RAND_896[1:0];
  _RAND_898 = {1{`RANDOM}};
  dataArray_18_11_cachedata_MPORT_en_pipe_0 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  dataArray_18_11_cachedata_MPORT_addr_pipe_0 = _RAND_899[1:0];
  _RAND_901 = {1{`RANDOM}};
  dataArray_18_12_cachedata_MPORT_en_pipe_0 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  dataArray_18_12_cachedata_MPORT_addr_pipe_0 = _RAND_902[1:0];
  _RAND_904 = {1{`RANDOM}};
  dataArray_18_13_cachedata_MPORT_en_pipe_0 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  dataArray_18_13_cachedata_MPORT_addr_pipe_0 = _RAND_905[1:0];
  _RAND_907 = {1{`RANDOM}};
  dataArray_18_14_cachedata_MPORT_en_pipe_0 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  dataArray_18_14_cachedata_MPORT_addr_pipe_0 = _RAND_908[1:0];
  _RAND_910 = {1{`RANDOM}};
  dataArray_18_15_cachedata_MPORT_en_pipe_0 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  dataArray_18_15_cachedata_MPORT_addr_pipe_0 = _RAND_911[1:0];
  _RAND_913 = {1{`RANDOM}};
  dataArray_19_0_cachedata_MPORT_en_pipe_0 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  dataArray_19_0_cachedata_MPORT_addr_pipe_0 = _RAND_914[1:0];
  _RAND_916 = {1{`RANDOM}};
  dataArray_19_1_cachedata_MPORT_en_pipe_0 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  dataArray_19_1_cachedata_MPORT_addr_pipe_0 = _RAND_917[1:0];
  _RAND_919 = {1{`RANDOM}};
  dataArray_19_2_cachedata_MPORT_en_pipe_0 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  dataArray_19_2_cachedata_MPORT_addr_pipe_0 = _RAND_920[1:0];
  _RAND_922 = {1{`RANDOM}};
  dataArray_19_3_cachedata_MPORT_en_pipe_0 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  dataArray_19_3_cachedata_MPORT_addr_pipe_0 = _RAND_923[1:0];
  _RAND_925 = {1{`RANDOM}};
  dataArray_19_4_cachedata_MPORT_en_pipe_0 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  dataArray_19_4_cachedata_MPORT_addr_pipe_0 = _RAND_926[1:0];
  _RAND_928 = {1{`RANDOM}};
  dataArray_19_5_cachedata_MPORT_en_pipe_0 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  dataArray_19_5_cachedata_MPORT_addr_pipe_0 = _RAND_929[1:0];
  _RAND_931 = {1{`RANDOM}};
  dataArray_19_6_cachedata_MPORT_en_pipe_0 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  dataArray_19_6_cachedata_MPORT_addr_pipe_0 = _RAND_932[1:0];
  _RAND_934 = {1{`RANDOM}};
  dataArray_19_7_cachedata_MPORT_en_pipe_0 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  dataArray_19_7_cachedata_MPORT_addr_pipe_0 = _RAND_935[1:0];
  _RAND_937 = {1{`RANDOM}};
  dataArray_19_8_cachedata_MPORT_en_pipe_0 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  dataArray_19_8_cachedata_MPORT_addr_pipe_0 = _RAND_938[1:0];
  _RAND_940 = {1{`RANDOM}};
  dataArray_19_9_cachedata_MPORT_en_pipe_0 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  dataArray_19_9_cachedata_MPORT_addr_pipe_0 = _RAND_941[1:0];
  _RAND_943 = {1{`RANDOM}};
  dataArray_19_10_cachedata_MPORT_en_pipe_0 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  dataArray_19_10_cachedata_MPORT_addr_pipe_0 = _RAND_944[1:0];
  _RAND_946 = {1{`RANDOM}};
  dataArray_19_11_cachedata_MPORT_en_pipe_0 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  dataArray_19_11_cachedata_MPORT_addr_pipe_0 = _RAND_947[1:0];
  _RAND_949 = {1{`RANDOM}};
  dataArray_19_12_cachedata_MPORT_en_pipe_0 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  dataArray_19_12_cachedata_MPORT_addr_pipe_0 = _RAND_950[1:0];
  _RAND_952 = {1{`RANDOM}};
  dataArray_19_13_cachedata_MPORT_en_pipe_0 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  dataArray_19_13_cachedata_MPORT_addr_pipe_0 = _RAND_953[1:0];
  _RAND_955 = {1{`RANDOM}};
  dataArray_19_14_cachedata_MPORT_en_pipe_0 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  dataArray_19_14_cachedata_MPORT_addr_pipe_0 = _RAND_956[1:0];
  _RAND_958 = {1{`RANDOM}};
  dataArray_19_15_cachedata_MPORT_en_pipe_0 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  dataArray_19_15_cachedata_MPORT_addr_pipe_0 = _RAND_959[1:0];
  _RAND_961 = {1{`RANDOM}};
  dataArray_20_0_cachedata_MPORT_en_pipe_0 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  dataArray_20_0_cachedata_MPORT_addr_pipe_0 = _RAND_962[1:0];
  _RAND_964 = {1{`RANDOM}};
  dataArray_20_1_cachedata_MPORT_en_pipe_0 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  dataArray_20_1_cachedata_MPORT_addr_pipe_0 = _RAND_965[1:0];
  _RAND_967 = {1{`RANDOM}};
  dataArray_20_2_cachedata_MPORT_en_pipe_0 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  dataArray_20_2_cachedata_MPORT_addr_pipe_0 = _RAND_968[1:0];
  _RAND_970 = {1{`RANDOM}};
  dataArray_20_3_cachedata_MPORT_en_pipe_0 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  dataArray_20_3_cachedata_MPORT_addr_pipe_0 = _RAND_971[1:0];
  _RAND_973 = {1{`RANDOM}};
  dataArray_20_4_cachedata_MPORT_en_pipe_0 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  dataArray_20_4_cachedata_MPORT_addr_pipe_0 = _RAND_974[1:0];
  _RAND_976 = {1{`RANDOM}};
  dataArray_20_5_cachedata_MPORT_en_pipe_0 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  dataArray_20_5_cachedata_MPORT_addr_pipe_0 = _RAND_977[1:0];
  _RAND_979 = {1{`RANDOM}};
  dataArray_20_6_cachedata_MPORT_en_pipe_0 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  dataArray_20_6_cachedata_MPORT_addr_pipe_0 = _RAND_980[1:0];
  _RAND_982 = {1{`RANDOM}};
  dataArray_20_7_cachedata_MPORT_en_pipe_0 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  dataArray_20_7_cachedata_MPORT_addr_pipe_0 = _RAND_983[1:0];
  _RAND_985 = {1{`RANDOM}};
  dataArray_20_8_cachedata_MPORT_en_pipe_0 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  dataArray_20_8_cachedata_MPORT_addr_pipe_0 = _RAND_986[1:0];
  _RAND_988 = {1{`RANDOM}};
  dataArray_20_9_cachedata_MPORT_en_pipe_0 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  dataArray_20_9_cachedata_MPORT_addr_pipe_0 = _RAND_989[1:0];
  _RAND_991 = {1{`RANDOM}};
  dataArray_20_10_cachedata_MPORT_en_pipe_0 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  dataArray_20_10_cachedata_MPORT_addr_pipe_0 = _RAND_992[1:0];
  _RAND_994 = {1{`RANDOM}};
  dataArray_20_11_cachedata_MPORT_en_pipe_0 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  dataArray_20_11_cachedata_MPORT_addr_pipe_0 = _RAND_995[1:0];
  _RAND_997 = {1{`RANDOM}};
  dataArray_20_12_cachedata_MPORT_en_pipe_0 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  dataArray_20_12_cachedata_MPORT_addr_pipe_0 = _RAND_998[1:0];
  _RAND_1000 = {1{`RANDOM}};
  dataArray_20_13_cachedata_MPORT_en_pipe_0 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  dataArray_20_13_cachedata_MPORT_addr_pipe_0 = _RAND_1001[1:0];
  _RAND_1003 = {1{`RANDOM}};
  dataArray_20_14_cachedata_MPORT_en_pipe_0 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  dataArray_20_14_cachedata_MPORT_addr_pipe_0 = _RAND_1004[1:0];
  _RAND_1006 = {1{`RANDOM}};
  dataArray_20_15_cachedata_MPORT_en_pipe_0 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  dataArray_20_15_cachedata_MPORT_addr_pipe_0 = _RAND_1007[1:0];
  _RAND_1009 = {1{`RANDOM}};
  dataArray_21_0_cachedata_MPORT_en_pipe_0 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  dataArray_21_0_cachedata_MPORT_addr_pipe_0 = _RAND_1010[1:0];
  _RAND_1012 = {1{`RANDOM}};
  dataArray_21_1_cachedata_MPORT_en_pipe_0 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  dataArray_21_1_cachedata_MPORT_addr_pipe_0 = _RAND_1013[1:0];
  _RAND_1015 = {1{`RANDOM}};
  dataArray_21_2_cachedata_MPORT_en_pipe_0 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  dataArray_21_2_cachedata_MPORT_addr_pipe_0 = _RAND_1016[1:0];
  _RAND_1018 = {1{`RANDOM}};
  dataArray_21_3_cachedata_MPORT_en_pipe_0 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  dataArray_21_3_cachedata_MPORT_addr_pipe_0 = _RAND_1019[1:0];
  _RAND_1021 = {1{`RANDOM}};
  dataArray_21_4_cachedata_MPORT_en_pipe_0 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  dataArray_21_4_cachedata_MPORT_addr_pipe_0 = _RAND_1022[1:0];
  _RAND_1024 = {1{`RANDOM}};
  dataArray_21_5_cachedata_MPORT_en_pipe_0 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  dataArray_21_5_cachedata_MPORT_addr_pipe_0 = _RAND_1025[1:0];
  _RAND_1027 = {1{`RANDOM}};
  dataArray_21_6_cachedata_MPORT_en_pipe_0 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  dataArray_21_6_cachedata_MPORT_addr_pipe_0 = _RAND_1028[1:0];
  _RAND_1030 = {1{`RANDOM}};
  dataArray_21_7_cachedata_MPORT_en_pipe_0 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  dataArray_21_7_cachedata_MPORT_addr_pipe_0 = _RAND_1031[1:0];
  _RAND_1033 = {1{`RANDOM}};
  dataArray_21_8_cachedata_MPORT_en_pipe_0 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  dataArray_21_8_cachedata_MPORT_addr_pipe_0 = _RAND_1034[1:0];
  _RAND_1036 = {1{`RANDOM}};
  dataArray_21_9_cachedata_MPORT_en_pipe_0 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  dataArray_21_9_cachedata_MPORT_addr_pipe_0 = _RAND_1037[1:0];
  _RAND_1039 = {1{`RANDOM}};
  dataArray_21_10_cachedata_MPORT_en_pipe_0 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  dataArray_21_10_cachedata_MPORT_addr_pipe_0 = _RAND_1040[1:0];
  _RAND_1042 = {1{`RANDOM}};
  dataArray_21_11_cachedata_MPORT_en_pipe_0 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  dataArray_21_11_cachedata_MPORT_addr_pipe_0 = _RAND_1043[1:0];
  _RAND_1045 = {1{`RANDOM}};
  dataArray_21_12_cachedata_MPORT_en_pipe_0 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  dataArray_21_12_cachedata_MPORT_addr_pipe_0 = _RAND_1046[1:0];
  _RAND_1048 = {1{`RANDOM}};
  dataArray_21_13_cachedata_MPORT_en_pipe_0 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  dataArray_21_13_cachedata_MPORT_addr_pipe_0 = _RAND_1049[1:0];
  _RAND_1051 = {1{`RANDOM}};
  dataArray_21_14_cachedata_MPORT_en_pipe_0 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  dataArray_21_14_cachedata_MPORT_addr_pipe_0 = _RAND_1052[1:0];
  _RAND_1054 = {1{`RANDOM}};
  dataArray_21_15_cachedata_MPORT_en_pipe_0 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  dataArray_21_15_cachedata_MPORT_addr_pipe_0 = _RAND_1055[1:0];
  _RAND_1057 = {1{`RANDOM}};
  dataArray_22_0_cachedata_MPORT_en_pipe_0 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  dataArray_22_0_cachedata_MPORT_addr_pipe_0 = _RAND_1058[1:0];
  _RAND_1060 = {1{`RANDOM}};
  dataArray_22_1_cachedata_MPORT_en_pipe_0 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  dataArray_22_1_cachedata_MPORT_addr_pipe_0 = _RAND_1061[1:0];
  _RAND_1063 = {1{`RANDOM}};
  dataArray_22_2_cachedata_MPORT_en_pipe_0 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  dataArray_22_2_cachedata_MPORT_addr_pipe_0 = _RAND_1064[1:0];
  _RAND_1066 = {1{`RANDOM}};
  dataArray_22_3_cachedata_MPORT_en_pipe_0 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  dataArray_22_3_cachedata_MPORT_addr_pipe_0 = _RAND_1067[1:0];
  _RAND_1069 = {1{`RANDOM}};
  dataArray_22_4_cachedata_MPORT_en_pipe_0 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  dataArray_22_4_cachedata_MPORT_addr_pipe_0 = _RAND_1070[1:0];
  _RAND_1072 = {1{`RANDOM}};
  dataArray_22_5_cachedata_MPORT_en_pipe_0 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  dataArray_22_5_cachedata_MPORT_addr_pipe_0 = _RAND_1073[1:0];
  _RAND_1075 = {1{`RANDOM}};
  dataArray_22_6_cachedata_MPORT_en_pipe_0 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  dataArray_22_6_cachedata_MPORT_addr_pipe_0 = _RAND_1076[1:0];
  _RAND_1078 = {1{`RANDOM}};
  dataArray_22_7_cachedata_MPORT_en_pipe_0 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  dataArray_22_7_cachedata_MPORT_addr_pipe_0 = _RAND_1079[1:0];
  _RAND_1081 = {1{`RANDOM}};
  dataArray_22_8_cachedata_MPORT_en_pipe_0 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  dataArray_22_8_cachedata_MPORT_addr_pipe_0 = _RAND_1082[1:0];
  _RAND_1084 = {1{`RANDOM}};
  dataArray_22_9_cachedata_MPORT_en_pipe_0 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  dataArray_22_9_cachedata_MPORT_addr_pipe_0 = _RAND_1085[1:0];
  _RAND_1087 = {1{`RANDOM}};
  dataArray_22_10_cachedata_MPORT_en_pipe_0 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  dataArray_22_10_cachedata_MPORT_addr_pipe_0 = _RAND_1088[1:0];
  _RAND_1090 = {1{`RANDOM}};
  dataArray_22_11_cachedata_MPORT_en_pipe_0 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  dataArray_22_11_cachedata_MPORT_addr_pipe_0 = _RAND_1091[1:0];
  _RAND_1093 = {1{`RANDOM}};
  dataArray_22_12_cachedata_MPORT_en_pipe_0 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  dataArray_22_12_cachedata_MPORT_addr_pipe_0 = _RAND_1094[1:0];
  _RAND_1096 = {1{`RANDOM}};
  dataArray_22_13_cachedata_MPORT_en_pipe_0 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  dataArray_22_13_cachedata_MPORT_addr_pipe_0 = _RAND_1097[1:0];
  _RAND_1099 = {1{`RANDOM}};
  dataArray_22_14_cachedata_MPORT_en_pipe_0 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  dataArray_22_14_cachedata_MPORT_addr_pipe_0 = _RAND_1100[1:0];
  _RAND_1102 = {1{`RANDOM}};
  dataArray_22_15_cachedata_MPORT_en_pipe_0 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  dataArray_22_15_cachedata_MPORT_addr_pipe_0 = _RAND_1103[1:0];
  _RAND_1105 = {1{`RANDOM}};
  dataArray_23_0_cachedata_MPORT_en_pipe_0 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  dataArray_23_0_cachedata_MPORT_addr_pipe_0 = _RAND_1106[1:0];
  _RAND_1108 = {1{`RANDOM}};
  dataArray_23_1_cachedata_MPORT_en_pipe_0 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  dataArray_23_1_cachedata_MPORT_addr_pipe_0 = _RAND_1109[1:0];
  _RAND_1111 = {1{`RANDOM}};
  dataArray_23_2_cachedata_MPORT_en_pipe_0 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  dataArray_23_2_cachedata_MPORT_addr_pipe_0 = _RAND_1112[1:0];
  _RAND_1114 = {1{`RANDOM}};
  dataArray_23_3_cachedata_MPORT_en_pipe_0 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  dataArray_23_3_cachedata_MPORT_addr_pipe_0 = _RAND_1115[1:0];
  _RAND_1117 = {1{`RANDOM}};
  dataArray_23_4_cachedata_MPORT_en_pipe_0 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  dataArray_23_4_cachedata_MPORT_addr_pipe_0 = _RAND_1118[1:0];
  _RAND_1120 = {1{`RANDOM}};
  dataArray_23_5_cachedata_MPORT_en_pipe_0 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  dataArray_23_5_cachedata_MPORT_addr_pipe_0 = _RAND_1121[1:0];
  _RAND_1123 = {1{`RANDOM}};
  dataArray_23_6_cachedata_MPORT_en_pipe_0 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  dataArray_23_6_cachedata_MPORT_addr_pipe_0 = _RAND_1124[1:0];
  _RAND_1126 = {1{`RANDOM}};
  dataArray_23_7_cachedata_MPORT_en_pipe_0 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  dataArray_23_7_cachedata_MPORT_addr_pipe_0 = _RAND_1127[1:0];
  _RAND_1129 = {1{`RANDOM}};
  dataArray_23_8_cachedata_MPORT_en_pipe_0 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  dataArray_23_8_cachedata_MPORT_addr_pipe_0 = _RAND_1130[1:0];
  _RAND_1132 = {1{`RANDOM}};
  dataArray_23_9_cachedata_MPORT_en_pipe_0 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  dataArray_23_9_cachedata_MPORT_addr_pipe_0 = _RAND_1133[1:0];
  _RAND_1135 = {1{`RANDOM}};
  dataArray_23_10_cachedata_MPORT_en_pipe_0 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  dataArray_23_10_cachedata_MPORT_addr_pipe_0 = _RAND_1136[1:0];
  _RAND_1138 = {1{`RANDOM}};
  dataArray_23_11_cachedata_MPORT_en_pipe_0 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  dataArray_23_11_cachedata_MPORT_addr_pipe_0 = _RAND_1139[1:0];
  _RAND_1141 = {1{`RANDOM}};
  dataArray_23_12_cachedata_MPORT_en_pipe_0 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  dataArray_23_12_cachedata_MPORT_addr_pipe_0 = _RAND_1142[1:0];
  _RAND_1144 = {1{`RANDOM}};
  dataArray_23_13_cachedata_MPORT_en_pipe_0 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  dataArray_23_13_cachedata_MPORT_addr_pipe_0 = _RAND_1145[1:0];
  _RAND_1147 = {1{`RANDOM}};
  dataArray_23_14_cachedata_MPORT_en_pipe_0 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  dataArray_23_14_cachedata_MPORT_addr_pipe_0 = _RAND_1148[1:0];
  _RAND_1150 = {1{`RANDOM}};
  dataArray_23_15_cachedata_MPORT_en_pipe_0 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  dataArray_23_15_cachedata_MPORT_addr_pipe_0 = _RAND_1151[1:0];
  _RAND_1153 = {1{`RANDOM}};
  dataArray_24_0_cachedata_MPORT_en_pipe_0 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  dataArray_24_0_cachedata_MPORT_addr_pipe_0 = _RAND_1154[1:0];
  _RAND_1156 = {1{`RANDOM}};
  dataArray_24_1_cachedata_MPORT_en_pipe_0 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  dataArray_24_1_cachedata_MPORT_addr_pipe_0 = _RAND_1157[1:0];
  _RAND_1159 = {1{`RANDOM}};
  dataArray_24_2_cachedata_MPORT_en_pipe_0 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  dataArray_24_2_cachedata_MPORT_addr_pipe_0 = _RAND_1160[1:0];
  _RAND_1162 = {1{`RANDOM}};
  dataArray_24_3_cachedata_MPORT_en_pipe_0 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  dataArray_24_3_cachedata_MPORT_addr_pipe_0 = _RAND_1163[1:0];
  _RAND_1165 = {1{`RANDOM}};
  dataArray_24_4_cachedata_MPORT_en_pipe_0 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  dataArray_24_4_cachedata_MPORT_addr_pipe_0 = _RAND_1166[1:0];
  _RAND_1168 = {1{`RANDOM}};
  dataArray_24_5_cachedata_MPORT_en_pipe_0 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  dataArray_24_5_cachedata_MPORT_addr_pipe_0 = _RAND_1169[1:0];
  _RAND_1171 = {1{`RANDOM}};
  dataArray_24_6_cachedata_MPORT_en_pipe_0 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  dataArray_24_6_cachedata_MPORT_addr_pipe_0 = _RAND_1172[1:0];
  _RAND_1174 = {1{`RANDOM}};
  dataArray_24_7_cachedata_MPORT_en_pipe_0 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  dataArray_24_7_cachedata_MPORT_addr_pipe_0 = _RAND_1175[1:0];
  _RAND_1177 = {1{`RANDOM}};
  dataArray_24_8_cachedata_MPORT_en_pipe_0 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  dataArray_24_8_cachedata_MPORT_addr_pipe_0 = _RAND_1178[1:0];
  _RAND_1180 = {1{`RANDOM}};
  dataArray_24_9_cachedata_MPORT_en_pipe_0 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  dataArray_24_9_cachedata_MPORT_addr_pipe_0 = _RAND_1181[1:0];
  _RAND_1183 = {1{`RANDOM}};
  dataArray_24_10_cachedata_MPORT_en_pipe_0 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  dataArray_24_10_cachedata_MPORT_addr_pipe_0 = _RAND_1184[1:0];
  _RAND_1186 = {1{`RANDOM}};
  dataArray_24_11_cachedata_MPORT_en_pipe_0 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  dataArray_24_11_cachedata_MPORT_addr_pipe_0 = _RAND_1187[1:0];
  _RAND_1189 = {1{`RANDOM}};
  dataArray_24_12_cachedata_MPORT_en_pipe_0 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  dataArray_24_12_cachedata_MPORT_addr_pipe_0 = _RAND_1190[1:0];
  _RAND_1192 = {1{`RANDOM}};
  dataArray_24_13_cachedata_MPORT_en_pipe_0 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  dataArray_24_13_cachedata_MPORT_addr_pipe_0 = _RAND_1193[1:0];
  _RAND_1195 = {1{`RANDOM}};
  dataArray_24_14_cachedata_MPORT_en_pipe_0 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  dataArray_24_14_cachedata_MPORT_addr_pipe_0 = _RAND_1196[1:0];
  _RAND_1198 = {1{`RANDOM}};
  dataArray_24_15_cachedata_MPORT_en_pipe_0 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  dataArray_24_15_cachedata_MPORT_addr_pipe_0 = _RAND_1199[1:0];
  _RAND_1201 = {1{`RANDOM}};
  dataArray_25_0_cachedata_MPORT_en_pipe_0 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  dataArray_25_0_cachedata_MPORT_addr_pipe_0 = _RAND_1202[1:0];
  _RAND_1204 = {1{`RANDOM}};
  dataArray_25_1_cachedata_MPORT_en_pipe_0 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  dataArray_25_1_cachedata_MPORT_addr_pipe_0 = _RAND_1205[1:0];
  _RAND_1207 = {1{`RANDOM}};
  dataArray_25_2_cachedata_MPORT_en_pipe_0 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  dataArray_25_2_cachedata_MPORT_addr_pipe_0 = _RAND_1208[1:0];
  _RAND_1210 = {1{`RANDOM}};
  dataArray_25_3_cachedata_MPORT_en_pipe_0 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  dataArray_25_3_cachedata_MPORT_addr_pipe_0 = _RAND_1211[1:0];
  _RAND_1213 = {1{`RANDOM}};
  dataArray_25_4_cachedata_MPORT_en_pipe_0 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  dataArray_25_4_cachedata_MPORT_addr_pipe_0 = _RAND_1214[1:0];
  _RAND_1216 = {1{`RANDOM}};
  dataArray_25_5_cachedata_MPORT_en_pipe_0 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  dataArray_25_5_cachedata_MPORT_addr_pipe_0 = _RAND_1217[1:0];
  _RAND_1219 = {1{`RANDOM}};
  dataArray_25_6_cachedata_MPORT_en_pipe_0 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  dataArray_25_6_cachedata_MPORT_addr_pipe_0 = _RAND_1220[1:0];
  _RAND_1222 = {1{`RANDOM}};
  dataArray_25_7_cachedata_MPORT_en_pipe_0 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  dataArray_25_7_cachedata_MPORT_addr_pipe_0 = _RAND_1223[1:0];
  _RAND_1225 = {1{`RANDOM}};
  dataArray_25_8_cachedata_MPORT_en_pipe_0 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  dataArray_25_8_cachedata_MPORT_addr_pipe_0 = _RAND_1226[1:0];
  _RAND_1228 = {1{`RANDOM}};
  dataArray_25_9_cachedata_MPORT_en_pipe_0 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  dataArray_25_9_cachedata_MPORT_addr_pipe_0 = _RAND_1229[1:0];
  _RAND_1231 = {1{`RANDOM}};
  dataArray_25_10_cachedata_MPORT_en_pipe_0 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  dataArray_25_10_cachedata_MPORT_addr_pipe_0 = _RAND_1232[1:0];
  _RAND_1234 = {1{`RANDOM}};
  dataArray_25_11_cachedata_MPORT_en_pipe_0 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  dataArray_25_11_cachedata_MPORT_addr_pipe_0 = _RAND_1235[1:0];
  _RAND_1237 = {1{`RANDOM}};
  dataArray_25_12_cachedata_MPORT_en_pipe_0 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  dataArray_25_12_cachedata_MPORT_addr_pipe_0 = _RAND_1238[1:0];
  _RAND_1240 = {1{`RANDOM}};
  dataArray_25_13_cachedata_MPORT_en_pipe_0 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  dataArray_25_13_cachedata_MPORT_addr_pipe_0 = _RAND_1241[1:0];
  _RAND_1243 = {1{`RANDOM}};
  dataArray_25_14_cachedata_MPORT_en_pipe_0 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  dataArray_25_14_cachedata_MPORT_addr_pipe_0 = _RAND_1244[1:0];
  _RAND_1246 = {1{`RANDOM}};
  dataArray_25_15_cachedata_MPORT_en_pipe_0 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  dataArray_25_15_cachedata_MPORT_addr_pipe_0 = _RAND_1247[1:0];
  _RAND_1249 = {1{`RANDOM}};
  dataArray_26_0_cachedata_MPORT_en_pipe_0 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  dataArray_26_0_cachedata_MPORT_addr_pipe_0 = _RAND_1250[1:0];
  _RAND_1252 = {1{`RANDOM}};
  dataArray_26_1_cachedata_MPORT_en_pipe_0 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  dataArray_26_1_cachedata_MPORT_addr_pipe_0 = _RAND_1253[1:0];
  _RAND_1255 = {1{`RANDOM}};
  dataArray_26_2_cachedata_MPORT_en_pipe_0 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  dataArray_26_2_cachedata_MPORT_addr_pipe_0 = _RAND_1256[1:0];
  _RAND_1258 = {1{`RANDOM}};
  dataArray_26_3_cachedata_MPORT_en_pipe_0 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  dataArray_26_3_cachedata_MPORT_addr_pipe_0 = _RAND_1259[1:0];
  _RAND_1261 = {1{`RANDOM}};
  dataArray_26_4_cachedata_MPORT_en_pipe_0 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  dataArray_26_4_cachedata_MPORT_addr_pipe_0 = _RAND_1262[1:0];
  _RAND_1264 = {1{`RANDOM}};
  dataArray_26_5_cachedata_MPORT_en_pipe_0 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  dataArray_26_5_cachedata_MPORT_addr_pipe_0 = _RAND_1265[1:0];
  _RAND_1267 = {1{`RANDOM}};
  dataArray_26_6_cachedata_MPORT_en_pipe_0 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  dataArray_26_6_cachedata_MPORT_addr_pipe_0 = _RAND_1268[1:0];
  _RAND_1270 = {1{`RANDOM}};
  dataArray_26_7_cachedata_MPORT_en_pipe_0 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  dataArray_26_7_cachedata_MPORT_addr_pipe_0 = _RAND_1271[1:0];
  _RAND_1273 = {1{`RANDOM}};
  dataArray_26_8_cachedata_MPORT_en_pipe_0 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  dataArray_26_8_cachedata_MPORT_addr_pipe_0 = _RAND_1274[1:0];
  _RAND_1276 = {1{`RANDOM}};
  dataArray_26_9_cachedata_MPORT_en_pipe_0 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  dataArray_26_9_cachedata_MPORT_addr_pipe_0 = _RAND_1277[1:0];
  _RAND_1279 = {1{`RANDOM}};
  dataArray_26_10_cachedata_MPORT_en_pipe_0 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  dataArray_26_10_cachedata_MPORT_addr_pipe_0 = _RAND_1280[1:0];
  _RAND_1282 = {1{`RANDOM}};
  dataArray_26_11_cachedata_MPORT_en_pipe_0 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  dataArray_26_11_cachedata_MPORT_addr_pipe_0 = _RAND_1283[1:0];
  _RAND_1285 = {1{`RANDOM}};
  dataArray_26_12_cachedata_MPORT_en_pipe_0 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  dataArray_26_12_cachedata_MPORT_addr_pipe_0 = _RAND_1286[1:0];
  _RAND_1288 = {1{`RANDOM}};
  dataArray_26_13_cachedata_MPORT_en_pipe_0 = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  dataArray_26_13_cachedata_MPORT_addr_pipe_0 = _RAND_1289[1:0];
  _RAND_1291 = {1{`RANDOM}};
  dataArray_26_14_cachedata_MPORT_en_pipe_0 = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  dataArray_26_14_cachedata_MPORT_addr_pipe_0 = _RAND_1292[1:0];
  _RAND_1294 = {1{`RANDOM}};
  dataArray_26_15_cachedata_MPORT_en_pipe_0 = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  dataArray_26_15_cachedata_MPORT_addr_pipe_0 = _RAND_1295[1:0];
  _RAND_1297 = {1{`RANDOM}};
  dataArray_27_0_cachedata_MPORT_en_pipe_0 = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  dataArray_27_0_cachedata_MPORT_addr_pipe_0 = _RAND_1298[1:0];
  _RAND_1300 = {1{`RANDOM}};
  dataArray_27_1_cachedata_MPORT_en_pipe_0 = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  dataArray_27_1_cachedata_MPORT_addr_pipe_0 = _RAND_1301[1:0];
  _RAND_1303 = {1{`RANDOM}};
  dataArray_27_2_cachedata_MPORT_en_pipe_0 = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  dataArray_27_2_cachedata_MPORT_addr_pipe_0 = _RAND_1304[1:0];
  _RAND_1306 = {1{`RANDOM}};
  dataArray_27_3_cachedata_MPORT_en_pipe_0 = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  dataArray_27_3_cachedata_MPORT_addr_pipe_0 = _RAND_1307[1:0];
  _RAND_1309 = {1{`RANDOM}};
  dataArray_27_4_cachedata_MPORT_en_pipe_0 = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  dataArray_27_4_cachedata_MPORT_addr_pipe_0 = _RAND_1310[1:0];
  _RAND_1312 = {1{`RANDOM}};
  dataArray_27_5_cachedata_MPORT_en_pipe_0 = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  dataArray_27_5_cachedata_MPORT_addr_pipe_0 = _RAND_1313[1:0];
  _RAND_1315 = {1{`RANDOM}};
  dataArray_27_6_cachedata_MPORT_en_pipe_0 = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  dataArray_27_6_cachedata_MPORT_addr_pipe_0 = _RAND_1316[1:0];
  _RAND_1318 = {1{`RANDOM}};
  dataArray_27_7_cachedata_MPORT_en_pipe_0 = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  dataArray_27_7_cachedata_MPORT_addr_pipe_0 = _RAND_1319[1:0];
  _RAND_1321 = {1{`RANDOM}};
  dataArray_27_8_cachedata_MPORT_en_pipe_0 = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  dataArray_27_8_cachedata_MPORT_addr_pipe_0 = _RAND_1322[1:0];
  _RAND_1324 = {1{`RANDOM}};
  dataArray_27_9_cachedata_MPORT_en_pipe_0 = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  dataArray_27_9_cachedata_MPORT_addr_pipe_0 = _RAND_1325[1:0];
  _RAND_1327 = {1{`RANDOM}};
  dataArray_27_10_cachedata_MPORT_en_pipe_0 = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  dataArray_27_10_cachedata_MPORT_addr_pipe_0 = _RAND_1328[1:0];
  _RAND_1330 = {1{`RANDOM}};
  dataArray_27_11_cachedata_MPORT_en_pipe_0 = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  dataArray_27_11_cachedata_MPORT_addr_pipe_0 = _RAND_1331[1:0];
  _RAND_1333 = {1{`RANDOM}};
  dataArray_27_12_cachedata_MPORT_en_pipe_0 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  dataArray_27_12_cachedata_MPORT_addr_pipe_0 = _RAND_1334[1:0];
  _RAND_1336 = {1{`RANDOM}};
  dataArray_27_13_cachedata_MPORT_en_pipe_0 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  dataArray_27_13_cachedata_MPORT_addr_pipe_0 = _RAND_1337[1:0];
  _RAND_1339 = {1{`RANDOM}};
  dataArray_27_14_cachedata_MPORT_en_pipe_0 = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  dataArray_27_14_cachedata_MPORT_addr_pipe_0 = _RAND_1340[1:0];
  _RAND_1342 = {1{`RANDOM}};
  dataArray_27_15_cachedata_MPORT_en_pipe_0 = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  dataArray_27_15_cachedata_MPORT_addr_pipe_0 = _RAND_1343[1:0];
  _RAND_1345 = {1{`RANDOM}};
  dataArray_28_0_cachedata_MPORT_en_pipe_0 = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  dataArray_28_0_cachedata_MPORT_addr_pipe_0 = _RAND_1346[1:0];
  _RAND_1348 = {1{`RANDOM}};
  dataArray_28_1_cachedata_MPORT_en_pipe_0 = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  dataArray_28_1_cachedata_MPORT_addr_pipe_0 = _RAND_1349[1:0];
  _RAND_1351 = {1{`RANDOM}};
  dataArray_28_2_cachedata_MPORT_en_pipe_0 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  dataArray_28_2_cachedata_MPORT_addr_pipe_0 = _RAND_1352[1:0];
  _RAND_1354 = {1{`RANDOM}};
  dataArray_28_3_cachedata_MPORT_en_pipe_0 = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  dataArray_28_3_cachedata_MPORT_addr_pipe_0 = _RAND_1355[1:0];
  _RAND_1357 = {1{`RANDOM}};
  dataArray_28_4_cachedata_MPORT_en_pipe_0 = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  dataArray_28_4_cachedata_MPORT_addr_pipe_0 = _RAND_1358[1:0];
  _RAND_1360 = {1{`RANDOM}};
  dataArray_28_5_cachedata_MPORT_en_pipe_0 = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  dataArray_28_5_cachedata_MPORT_addr_pipe_0 = _RAND_1361[1:0];
  _RAND_1363 = {1{`RANDOM}};
  dataArray_28_6_cachedata_MPORT_en_pipe_0 = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  dataArray_28_6_cachedata_MPORT_addr_pipe_0 = _RAND_1364[1:0];
  _RAND_1366 = {1{`RANDOM}};
  dataArray_28_7_cachedata_MPORT_en_pipe_0 = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  dataArray_28_7_cachedata_MPORT_addr_pipe_0 = _RAND_1367[1:0];
  _RAND_1369 = {1{`RANDOM}};
  dataArray_28_8_cachedata_MPORT_en_pipe_0 = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  dataArray_28_8_cachedata_MPORT_addr_pipe_0 = _RAND_1370[1:0];
  _RAND_1372 = {1{`RANDOM}};
  dataArray_28_9_cachedata_MPORT_en_pipe_0 = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  dataArray_28_9_cachedata_MPORT_addr_pipe_0 = _RAND_1373[1:0];
  _RAND_1375 = {1{`RANDOM}};
  dataArray_28_10_cachedata_MPORT_en_pipe_0 = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  dataArray_28_10_cachedata_MPORT_addr_pipe_0 = _RAND_1376[1:0];
  _RAND_1378 = {1{`RANDOM}};
  dataArray_28_11_cachedata_MPORT_en_pipe_0 = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  dataArray_28_11_cachedata_MPORT_addr_pipe_0 = _RAND_1379[1:0];
  _RAND_1381 = {1{`RANDOM}};
  dataArray_28_12_cachedata_MPORT_en_pipe_0 = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  dataArray_28_12_cachedata_MPORT_addr_pipe_0 = _RAND_1382[1:0];
  _RAND_1384 = {1{`RANDOM}};
  dataArray_28_13_cachedata_MPORT_en_pipe_0 = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  dataArray_28_13_cachedata_MPORT_addr_pipe_0 = _RAND_1385[1:0];
  _RAND_1387 = {1{`RANDOM}};
  dataArray_28_14_cachedata_MPORT_en_pipe_0 = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  dataArray_28_14_cachedata_MPORT_addr_pipe_0 = _RAND_1388[1:0];
  _RAND_1390 = {1{`RANDOM}};
  dataArray_28_15_cachedata_MPORT_en_pipe_0 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  dataArray_28_15_cachedata_MPORT_addr_pipe_0 = _RAND_1391[1:0];
  _RAND_1393 = {1{`RANDOM}};
  dataArray_29_0_cachedata_MPORT_en_pipe_0 = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  dataArray_29_0_cachedata_MPORT_addr_pipe_0 = _RAND_1394[1:0];
  _RAND_1396 = {1{`RANDOM}};
  dataArray_29_1_cachedata_MPORT_en_pipe_0 = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  dataArray_29_1_cachedata_MPORT_addr_pipe_0 = _RAND_1397[1:0];
  _RAND_1399 = {1{`RANDOM}};
  dataArray_29_2_cachedata_MPORT_en_pipe_0 = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  dataArray_29_2_cachedata_MPORT_addr_pipe_0 = _RAND_1400[1:0];
  _RAND_1402 = {1{`RANDOM}};
  dataArray_29_3_cachedata_MPORT_en_pipe_0 = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  dataArray_29_3_cachedata_MPORT_addr_pipe_0 = _RAND_1403[1:0];
  _RAND_1405 = {1{`RANDOM}};
  dataArray_29_4_cachedata_MPORT_en_pipe_0 = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  dataArray_29_4_cachedata_MPORT_addr_pipe_0 = _RAND_1406[1:0];
  _RAND_1408 = {1{`RANDOM}};
  dataArray_29_5_cachedata_MPORT_en_pipe_0 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  dataArray_29_5_cachedata_MPORT_addr_pipe_0 = _RAND_1409[1:0];
  _RAND_1411 = {1{`RANDOM}};
  dataArray_29_6_cachedata_MPORT_en_pipe_0 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  dataArray_29_6_cachedata_MPORT_addr_pipe_0 = _RAND_1412[1:0];
  _RAND_1414 = {1{`RANDOM}};
  dataArray_29_7_cachedata_MPORT_en_pipe_0 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  dataArray_29_7_cachedata_MPORT_addr_pipe_0 = _RAND_1415[1:0];
  _RAND_1417 = {1{`RANDOM}};
  dataArray_29_8_cachedata_MPORT_en_pipe_0 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  dataArray_29_8_cachedata_MPORT_addr_pipe_0 = _RAND_1418[1:0];
  _RAND_1420 = {1{`RANDOM}};
  dataArray_29_9_cachedata_MPORT_en_pipe_0 = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  dataArray_29_9_cachedata_MPORT_addr_pipe_0 = _RAND_1421[1:0];
  _RAND_1423 = {1{`RANDOM}};
  dataArray_29_10_cachedata_MPORT_en_pipe_0 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  dataArray_29_10_cachedata_MPORT_addr_pipe_0 = _RAND_1424[1:0];
  _RAND_1426 = {1{`RANDOM}};
  dataArray_29_11_cachedata_MPORT_en_pipe_0 = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  dataArray_29_11_cachedata_MPORT_addr_pipe_0 = _RAND_1427[1:0];
  _RAND_1429 = {1{`RANDOM}};
  dataArray_29_12_cachedata_MPORT_en_pipe_0 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  dataArray_29_12_cachedata_MPORT_addr_pipe_0 = _RAND_1430[1:0];
  _RAND_1432 = {1{`RANDOM}};
  dataArray_29_13_cachedata_MPORT_en_pipe_0 = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  dataArray_29_13_cachedata_MPORT_addr_pipe_0 = _RAND_1433[1:0];
  _RAND_1435 = {1{`RANDOM}};
  dataArray_29_14_cachedata_MPORT_en_pipe_0 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  dataArray_29_14_cachedata_MPORT_addr_pipe_0 = _RAND_1436[1:0];
  _RAND_1438 = {1{`RANDOM}};
  dataArray_29_15_cachedata_MPORT_en_pipe_0 = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  dataArray_29_15_cachedata_MPORT_addr_pipe_0 = _RAND_1439[1:0];
  _RAND_1441 = {1{`RANDOM}};
  dataArray_30_0_cachedata_MPORT_en_pipe_0 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  dataArray_30_0_cachedata_MPORT_addr_pipe_0 = _RAND_1442[1:0];
  _RAND_1444 = {1{`RANDOM}};
  dataArray_30_1_cachedata_MPORT_en_pipe_0 = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  dataArray_30_1_cachedata_MPORT_addr_pipe_0 = _RAND_1445[1:0];
  _RAND_1447 = {1{`RANDOM}};
  dataArray_30_2_cachedata_MPORT_en_pipe_0 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  dataArray_30_2_cachedata_MPORT_addr_pipe_0 = _RAND_1448[1:0];
  _RAND_1450 = {1{`RANDOM}};
  dataArray_30_3_cachedata_MPORT_en_pipe_0 = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  dataArray_30_3_cachedata_MPORT_addr_pipe_0 = _RAND_1451[1:0];
  _RAND_1453 = {1{`RANDOM}};
  dataArray_30_4_cachedata_MPORT_en_pipe_0 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  dataArray_30_4_cachedata_MPORT_addr_pipe_0 = _RAND_1454[1:0];
  _RAND_1456 = {1{`RANDOM}};
  dataArray_30_5_cachedata_MPORT_en_pipe_0 = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  dataArray_30_5_cachedata_MPORT_addr_pipe_0 = _RAND_1457[1:0];
  _RAND_1459 = {1{`RANDOM}};
  dataArray_30_6_cachedata_MPORT_en_pipe_0 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  dataArray_30_6_cachedata_MPORT_addr_pipe_0 = _RAND_1460[1:0];
  _RAND_1462 = {1{`RANDOM}};
  dataArray_30_7_cachedata_MPORT_en_pipe_0 = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  dataArray_30_7_cachedata_MPORT_addr_pipe_0 = _RAND_1463[1:0];
  _RAND_1465 = {1{`RANDOM}};
  dataArray_30_8_cachedata_MPORT_en_pipe_0 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  dataArray_30_8_cachedata_MPORT_addr_pipe_0 = _RAND_1466[1:0];
  _RAND_1468 = {1{`RANDOM}};
  dataArray_30_9_cachedata_MPORT_en_pipe_0 = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  dataArray_30_9_cachedata_MPORT_addr_pipe_0 = _RAND_1469[1:0];
  _RAND_1471 = {1{`RANDOM}};
  dataArray_30_10_cachedata_MPORT_en_pipe_0 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  dataArray_30_10_cachedata_MPORT_addr_pipe_0 = _RAND_1472[1:0];
  _RAND_1474 = {1{`RANDOM}};
  dataArray_30_11_cachedata_MPORT_en_pipe_0 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  dataArray_30_11_cachedata_MPORT_addr_pipe_0 = _RAND_1475[1:0];
  _RAND_1477 = {1{`RANDOM}};
  dataArray_30_12_cachedata_MPORT_en_pipe_0 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  dataArray_30_12_cachedata_MPORT_addr_pipe_0 = _RAND_1478[1:0];
  _RAND_1480 = {1{`RANDOM}};
  dataArray_30_13_cachedata_MPORT_en_pipe_0 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  dataArray_30_13_cachedata_MPORT_addr_pipe_0 = _RAND_1481[1:0];
  _RAND_1483 = {1{`RANDOM}};
  dataArray_30_14_cachedata_MPORT_en_pipe_0 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  dataArray_30_14_cachedata_MPORT_addr_pipe_0 = _RAND_1484[1:0];
  _RAND_1486 = {1{`RANDOM}};
  dataArray_30_15_cachedata_MPORT_en_pipe_0 = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  dataArray_30_15_cachedata_MPORT_addr_pipe_0 = _RAND_1487[1:0];
  _RAND_1489 = {1{`RANDOM}};
  dataArray_31_0_cachedata_MPORT_en_pipe_0 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  dataArray_31_0_cachedata_MPORT_addr_pipe_0 = _RAND_1490[1:0];
  _RAND_1492 = {1{`RANDOM}};
  dataArray_31_1_cachedata_MPORT_en_pipe_0 = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  dataArray_31_1_cachedata_MPORT_addr_pipe_0 = _RAND_1493[1:0];
  _RAND_1495 = {1{`RANDOM}};
  dataArray_31_2_cachedata_MPORT_en_pipe_0 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  dataArray_31_2_cachedata_MPORT_addr_pipe_0 = _RAND_1496[1:0];
  _RAND_1498 = {1{`RANDOM}};
  dataArray_31_3_cachedata_MPORT_en_pipe_0 = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  dataArray_31_3_cachedata_MPORT_addr_pipe_0 = _RAND_1499[1:0];
  _RAND_1501 = {1{`RANDOM}};
  dataArray_31_4_cachedata_MPORT_en_pipe_0 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  dataArray_31_4_cachedata_MPORT_addr_pipe_0 = _RAND_1502[1:0];
  _RAND_1504 = {1{`RANDOM}};
  dataArray_31_5_cachedata_MPORT_en_pipe_0 = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  dataArray_31_5_cachedata_MPORT_addr_pipe_0 = _RAND_1505[1:0];
  _RAND_1507 = {1{`RANDOM}};
  dataArray_31_6_cachedata_MPORT_en_pipe_0 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  dataArray_31_6_cachedata_MPORT_addr_pipe_0 = _RAND_1508[1:0];
  _RAND_1510 = {1{`RANDOM}};
  dataArray_31_7_cachedata_MPORT_en_pipe_0 = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  dataArray_31_7_cachedata_MPORT_addr_pipe_0 = _RAND_1511[1:0];
  _RAND_1513 = {1{`RANDOM}};
  dataArray_31_8_cachedata_MPORT_en_pipe_0 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  dataArray_31_8_cachedata_MPORT_addr_pipe_0 = _RAND_1514[1:0];
  _RAND_1516 = {1{`RANDOM}};
  dataArray_31_9_cachedata_MPORT_en_pipe_0 = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  dataArray_31_9_cachedata_MPORT_addr_pipe_0 = _RAND_1517[1:0];
  _RAND_1519 = {1{`RANDOM}};
  dataArray_31_10_cachedata_MPORT_en_pipe_0 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  dataArray_31_10_cachedata_MPORT_addr_pipe_0 = _RAND_1520[1:0];
  _RAND_1522 = {1{`RANDOM}};
  dataArray_31_11_cachedata_MPORT_en_pipe_0 = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  dataArray_31_11_cachedata_MPORT_addr_pipe_0 = _RAND_1523[1:0];
  _RAND_1525 = {1{`RANDOM}};
  dataArray_31_12_cachedata_MPORT_en_pipe_0 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  dataArray_31_12_cachedata_MPORT_addr_pipe_0 = _RAND_1526[1:0];
  _RAND_1528 = {1{`RANDOM}};
  dataArray_31_13_cachedata_MPORT_en_pipe_0 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  dataArray_31_13_cachedata_MPORT_addr_pipe_0 = _RAND_1529[1:0];
  _RAND_1531 = {1{`RANDOM}};
  dataArray_31_14_cachedata_MPORT_en_pipe_0 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  dataArray_31_14_cachedata_MPORT_addr_pipe_0 = _RAND_1532[1:0];
  _RAND_1534 = {1{`RANDOM}};
  dataArray_31_15_cachedata_MPORT_en_pipe_0 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  dataArray_31_15_cachedata_MPORT_addr_pipe_0 = _RAND_1535[1:0];
  _RAND_1537 = {1{`RANDOM}};
  dataArray_32_0_cachedata_MPORT_en_pipe_0 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  dataArray_32_0_cachedata_MPORT_addr_pipe_0 = _RAND_1538[1:0];
  _RAND_1540 = {1{`RANDOM}};
  dataArray_32_1_cachedata_MPORT_en_pipe_0 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  dataArray_32_1_cachedata_MPORT_addr_pipe_0 = _RAND_1541[1:0];
  _RAND_1543 = {1{`RANDOM}};
  dataArray_32_2_cachedata_MPORT_en_pipe_0 = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  dataArray_32_2_cachedata_MPORT_addr_pipe_0 = _RAND_1544[1:0];
  _RAND_1546 = {1{`RANDOM}};
  dataArray_32_3_cachedata_MPORT_en_pipe_0 = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  dataArray_32_3_cachedata_MPORT_addr_pipe_0 = _RAND_1547[1:0];
  _RAND_1549 = {1{`RANDOM}};
  dataArray_32_4_cachedata_MPORT_en_pipe_0 = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  dataArray_32_4_cachedata_MPORT_addr_pipe_0 = _RAND_1550[1:0];
  _RAND_1552 = {1{`RANDOM}};
  dataArray_32_5_cachedata_MPORT_en_pipe_0 = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  dataArray_32_5_cachedata_MPORT_addr_pipe_0 = _RAND_1553[1:0];
  _RAND_1555 = {1{`RANDOM}};
  dataArray_32_6_cachedata_MPORT_en_pipe_0 = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  dataArray_32_6_cachedata_MPORT_addr_pipe_0 = _RAND_1556[1:0];
  _RAND_1558 = {1{`RANDOM}};
  dataArray_32_7_cachedata_MPORT_en_pipe_0 = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  dataArray_32_7_cachedata_MPORT_addr_pipe_0 = _RAND_1559[1:0];
  _RAND_1561 = {1{`RANDOM}};
  dataArray_32_8_cachedata_MPORT_en_pipe_0 = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  dataArray_32_8_cachedata_MPORT_addr_pipe_0 = _RAND_1562[1:0];
  _RAND_1564 = {1{`RANDOM}};
  dataArray_32_9_cachedata_MPORT_en_pipe_0 = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  dataArray_32_9_cachedata_MPORT_addr_pipe_0 = _RAND_1565[1:0];
  _RAND_1567 = {1{`RANDOM}};
  dataArray_32_10_cachedata_MPORT_en_pipe_0 = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  dataArray_32_10_cachedata_MPORT_addr_pipe_0 = _RAND_1568[1:0];
  _RAND_1570 = {1{`RANDOM}};
  dataArray_32_11_cachedata_MPORT_en_pipe_0 = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  dataArray_32_11_cachedata_MPORT_addr_pipe_0 = _RAND_1571[1:0];
  _RAND_1573 = {1{`RANDOM}};
  dataArray_32_12_cachedata_MPORT_en_pipe_0 = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  dataArray_32_12_cachedata_MPORT_addr_pipe_0 = _RAND_1574[1:0];
  _RAND_1576 = {1{`RANDOM}};
  dataArray_32_13_cachedata_MPORT_en_pipe_0 = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  dataArray_32_13_cachedata_MPORT_addr_pipe_0 = _RAND_1577[1:0];
  _RAND_1579 = {1{`RANDOM}};
  dataArray_32_14_cachedata_MPORT_en_pipe_0 = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  dataArray_32_14_cachedata_MPORT_addr_pipe_0 = _RAND_1580[1:0];
  _RAND_1582 = {1{`RANDOM}};
  dataArray_32_15_cachedata_MPORT_en_pipe_0 = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  dataArray_32_15_cachedata_MPORT_addr_pipe_0 = _RAND_1583[1:0];
  _RAND_1585 = {1{`RANDOM}};
  dataArray_33_0_cachedata_MPORT_en_pipe_0 = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  dataArray_33_0_cachedata_MPORT_addr_pipe_0 = _RAND_1586[1:0];
  _RAND_1588 = {1{`RANDOM}};
  dataArray_33_1_cachedata_MPORT_en_pipe_0 = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  dataArray_33_1_cachedata_MPORT_addr_pipe_0 = _RAND_1589[1:0];
  _RAND_1591 = {1{`RANDOM}};
  dataArray_33_2_cachedata_MPORT_en_pipe_0 = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  dataArray_33_2_cachedata_MPORT_addr_pipe_0 = _RAND_1592[1:0];
  _RAND_1594 = {1{`RANDOM}};
  dataArray_33_3_cachedata_MPORT_en_pipe_0 = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  dataArray_33_3_cachedata_MPORT_addr_pipe_0 = _RAND_1595[1:0];
  _RAND_1597 = {1{`RANDOM}};
  dataArray_33_4_cachedata_MPORT_en_pipe_0 = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  dataArray_33_4_cachedata_MPORT_addr_pipe_0 = _RAND_1598[1:0];
  _RAND_1600 = {1{`RANDOM}};
  dataArray_33_5_cachedata_MPORT_en_pipe_0 = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  dataArray_33_5_cachedata_MPORT_addr_pipe_0 = _RAND_1601[1:0];
  _RAND_1603 = {1{`RANDOM}};
  dataArray_33_6_cachedata_MPORT_en_pipe_0 = _RAND_1603[0:0];
  _RAND_1604 = {1{`RANDOM}};
  dataArray_33_6_cachedata_MPORT_addr_pipe_0 = _RAND_1604[1:0];
  _RAND_1606 = {1{`RANDOM}};
  dataArray_33_7_cachedata_MPORT_en_pipe_0 = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  dataArray_33_7_cachedata_MPORT_addr_pipe_0 = _RAND_1607[1:0];
  _RAND_1609 = {1{`RANDOM}};
  dataArray_33_8_cachedata_MPORT_en_pipe_0 = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  dataArray_33_8_cachedata_MPORT_addr_pipe_0 = _RAND_1610[1:0];
  _RAND_1612 = {1{`RANDOM}};
  dataArray_33_9_cachedata_MPORT_en_pipe_0 = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  dataArray_33_9_cachedata_MPORT_addr_pipe_0 = _RAND_1613[1:0];
  _RAND_1615 = {1{`RANDOM}};
  dataArray_33_10_cachedata_MPORT_en_pipe_0 = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  dataArray_33_10_cachedata_MPORT_addr_pipe_0 = _RAND_1616[1:0];
  _RAND_1618 = {1{`RANDOM}};
  dataArray_33_11_cachedata_MPORT_en_pipe_0 = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  dataArray_33_11_cachedata_MPORT_addr_pipe_0 = _RAND_1619[1:0];
  _RAND_1621 = {1{`RANDOM}};
  dataArray_33_12_cachedata_MPORT_en_pipe_0 = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  dataArray_33_12_cachedata_MPORT_addr_pipe_0 = _RAND_1622[1:0];
  _RAND_1624 = {1{`RANDOM}};
  dataArray_33_13_cachedata_MPORT_en_pipe_0 = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  dataArray_33_13_cachedata_MPORT_addr_pipe_0 = _RAND_1625[1:0];
  _RAND_1627 = {1{`RANDOM}};
  dataArray_33_14_cachedata_MPORT_en_pipe_0 = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  dataArray_33_14_cachedata_MPORT_addr_pipe_0 = _RAND_1628[1:0];
  _RAND_1630 = {1{`RANDOM}};
  dataArray_33_15_cachedata_MPORT_en_pipe_0 = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  dataArray_33_15_cachedata_MPORT_addr_pipe_0 = _RAND_1631[1:0];
  _RAND_1633 = {1{`RANDOM}};
  dataArray_34_0_cachedata_MPORT_en_pipe_0 = _RAND_1633[0:0];
  _RAND_1634 = {1{`RANDOM}};
  dataArray_34_0_cachedata_MPORT_addr_pipe_0 = _RAND_1634[1:0];
  _RAND_1636 = {1{`RANDOM}};
  dataArray_34_1_cachedata_MPORT_en_pipe_0 = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  dataArray_34_1_cachedata_MPORT_addr_pipe_0 = _RAND_1637[1:0];
  _RAND_1639 = {1{`RANDOM}};
  dataArray_34_2_cachedata_MPORT_en_pipe_0 = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  dataArray_34_2_cachedata_MPORT_addr_pipe_0 = _RAND_1640[1:0];
  _RAND_1642 = {1{`RANDOM}};
  dataArray_34_3_cachedata_MPORT_en_pipe_0 = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  dataArray_34_3_cachedata_MPORT_addr_pipe_0 = _RAND_1643[1:0];
  _RAND_1645 = {1{`RANDOM}};
  dataArray_34_4_cachedata_MPORT_en_pipe_0 = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  dataArray_34_4_cachedata_MPORT_addr_pipe_0 = _RAND_1646[1:0];
  _RAND_1648 = {1{`RANDOM}};
  dataArray_34_5_cachedata_MPORT_en_pipe_0 = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  dataArray_34_5_cachedata_MPORT_addr_pipe_0 = _RAND_1649[1:0];
  _RAND_1651 = {1{`RANDOM}};
  dataArray_34_6_cachedata_MPORT_en_pipe_0 = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  dataArray_34_6_cachedata_MPORT_addr_pipe_0 = _RAND_1652[1:0];
  _RAND_1654 = {1{`RANDOM}};
  dataArray_34_7_cachedata_MPORT_en_pipe_0 = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  dataArray_34_7_cachedata_MPORT_addr_pipe_0 = _RAND_1655[1:0];
  _RAND_1657 = {1{`RANDOM}};
  dataArray_34_8_cachedata_MPORT_en_pipe_0 = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  dataArray_34_8_cachedata_MPORT_addr_pipe_0 = _RAND_1658[1:0];
  _RAND_1660 = {1{`RANDOM}};
  dataArray_34_9_cachedata_MPORT_en_pipe_0 = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  dataArray_34_9_cachedata_MPORT_addr_pipe_0 = _RAND_1661[1:0];
  _RAND_1663 = {1{`RANDOM}};
  dataArray_34_10_cachedata_MPORT_en_pipe_0 = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  dataArray_34_10_cachedata_MPORT_addr_pipe_0 = _RAND_1664[1:0];
  _RAND_1666 = {1{`RANDOM}};
  dataArray_34_11_cachedata_MPORT_en_pipe_0 = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  dataArray_34_11_cachedata_MPORT_addr_pipe_0 = _RAND_1667[1:0];
  _RAND_1669 = {1{`RANDOM}};
  dataArray_34_12_cachedata_MPORT_en_pipe_0 = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  dataArray_34_12_cachedata_MPORT_addr_pipe_0 = _RAND_1670[1:0];
  _RAND_1672 = {1{`RANDOM}};
  dataArray_34_13_cachedata_MPORT_en_pipe_0 = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  dataArray_34_13_cachedata_MPORT_addr_pipe_0 = _RAND_1673[1:0];
  _RAND_1675 = {1{`RANDOM}};
  dataArray_34_14_cachedata_MPORT_en_pipe_0 = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  dataArray_34_14_cachedata_MPORT_addr_pipe_0 = _RAND_1676[1:0];
  _RAND_1678 = {1{`RANDOM}};
  dataArray_34_15_cachedata_MPORT_en_pipe_0 = _RAND_1678[0:0];
  _RAND_1679 = {1{`RANDOM}};
  dataArray_34_15_cachedata_MPORT_addr_pipe_0 = _RAND_1679[1:0];
  _RAND_1681 = {1{`RANDOM}};
  dataArray_35_0_cachedata_MPORT_en_pipe_0 = _RAND_1681[0:0];
  _RAND_1682 = {1{`RANDOM}};
  dataArray_35_0_cachedata_MPORT_addr_pipe_0 = _RAND_1682[1:0];
  _RAND_1684 = {1{`RANDOM}};
  dataArray_35_1_cachedata_MPORT_en_pipe_0 = _RAND_1684[0:0];
  _RAND_1685 = {1{`RANDOM}};
  dataArray_35_1_cachedata_MPORT_addr_pipe_0 = _RAND_1685[1:0];
  _RAND_1687 = {1{`RANDOM}};
  dataArray_35_2_cachedata_MPORT_en_pipe_0 = _RAND_1687[0:0];
  _RAND_1688 = {1{`RANDOM}};
  dataArray_35_2_cachedata_MPORT_addr_pipe_0 = _RAND_1688[1:0];
  _RAND_1690 = {1{`RANDOM}};
  dataArray_35_3_cachedata_MPORT_en_pipe_0 = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  dataArray_35_3_cachedata_MPORT_addr_pipe_0 = _RAND_1691[1:0];
  _RAND_1693 = {1{`RANDOM}};
  dataArray_35_4_cachedata_MPORT_en_pipe_0 = _RAND_1693[0:0];
  _RAND_1694 = {1{`RANDOM}};
  dataArray_35_4_cachedata_MPORT_addr_pipe_0 = _RAND_1694[1:0];
  _RAND_1696 = {1{`RANDOM}};
  dataArray_35_5_cachedata_MPORT_en_pipe_0 = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  dataArray_35_5_cachedata_MPORT_addr_pipe_0 = _RAND_1697[1:0];
  _RAND_1699 = {1{`RANDOM}};
  dataArray_35_6_cachedata_MPORT_en_pipe_0 = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  dataArray_35_6_cachedata_MPORT_addr_pipe_0 = _RAND_1700[1:0];
  _RAND_1702 = {1{`RANDOM}};
  dataArray_35_7_cachedata_MPORT_en_pipe_0 = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  dataArray_35_7_cachedata_MPORT_addr_pipe_0 = _RAND_1703[1:0];
  _RAND_1705 = {1{`RANDOM}};
  dataArray_35_8_cachedata_MPORT_en_pipe_0 = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  dataArray_35_8_cachedata_MPORT_addr_pipe_0 = _RAND_1706[1:0];
  _RAND_1708 = {1{`RANDOM}};
  dataArray_35_9_cachedata_MPORT_en_pipe_0 = _RAND_1708[0:0];
  _RAND_1709 = {1{`RANDOM}};
  dataArray_35_9_cachedata_MPORT_addr_pipe_0 = _RAND_1709[1:0];
  _RAND_1711 = {1{`RANDOM}};
  dataArray_35_10_cachedata_MPORT_en_pipe_0 = _RAND_1711[0:0];
  _RAND_1712 = {1{`RANDOM}};
  dataArray_35_10_cachedata_MPORT_addr_pipe_0 = _RAND_1712[1:0];
  _RAND_1714 = {1{`RANDOM}};
  dataArray_35_11_cachedata_MPORT_en_pipe_0 = _RAND_1714[0:0];
  _RAND_1715 = {1{`RANDOM}};
  dataArray_35_11_cachedata_MPORT_addr_pipe_0 = _RAND_1715[1:0];
  _RAND_1717 = {1{`RANDOM}};
  dataArray_35_12_cachedata_MPORT_en_pipe_0 = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  dataArray_35_12_cachedata_MPORT_addr_pipe_0 = _RAND_1718[1:0];
  _RAND_1720 = {1{`RANDOM}};
  dataArray_35_13_cachedata_MPORT_en_pipe_0 = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  dataArray_35_13_cachedata_MPORT_addr_pipe_0 = _RAND_1721[1:0];
  _RAND_1723 = {1{`RANDOM}};
  dataArray_35_14_cachedata_MPORT_en_pipe_0 = _RAND_1723[0:0];
  _RAND_1724 = {1{`RANDOM}};
  dataArray_35_14_cachedata_MPORT_addr_pipe_0 = _RAND_1724[1:0];
  _RAND_1726 = {1{`RANDOM}};
  dataArray_35_15_cachedata_MPORT_en_pipe_0 = _RAND_1726[0:0];
  _RAND_1727 = {1{`RANDOM}};
  dataArray_35_15_cachedata_MPORT_addr_pipe_0 = _RAND_1727[1:0];
  _RAND_1729 = {1{`RANDOM}};
  dataArray_36_0_cachedata_MPORT_en_pipe_0 = _RAND_1729[0:0];
  _RAND_1730 = {1{`RANDOM}};
  dataArray_36_0_cachedata_MPORT_addr_pipe_0 = _RAND_1730[1:0];
  _RAND_1732 = {1{`RANDOM}};
  dataArray_36_1_cachedata_MPORT_en_pipe_0 = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  dataArray_36_1_cachedata_MPORT_addr_pipe_0 = _RAND_1733[1:0];
  _RAND_1735 = {1{`RANDOM}};
  dataArray_36_2_cachedata_MPORT_en_pipe_0 = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  dataArray_36_2_cachedata_MPORT_addr_pipe_0 = _RAND_1736[1:0];
  _RAND_1738 = {1{`RANDOM}};
  dataArray_36_3_cachedata_MPORT_en_pipe_0 = _RAND_1738[0:0];
  _RAND_1739 = {1{`RANDOM}};
  dataArray_36_3_cachedata_MPORT_addr_pipe_0 = _RAND_1739[1:0];
  _RAND_1741 = {1{`RANDOM}};
  dataArray_36_4_cachedata_MPORT_en_pipe_0 = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  dataArray_36_4_cachedata_MPORT_addr_pipe_0 = _RAND_1742[1:0];
  _RAND_1744 = {1{`RANDOM}};
  dataArray_36_5_cachedata_MPORT_en_pipe_0 = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  dataArray_36_5_cachedata_MPORT_addr_pipe_0 = _RAND_1745[1:0];
  _RAND_1747 = {1{`RANDOM}};
  dataArray_36_6_cachedata_MPORT_en_pipe_0 = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  dataArray_36_6_cachedata_MPORT_addr_pipe_0 = _RAND_1748[1:0];
  _RAND_1750 = {1{`RANDOM}};
  dataArray_36_7_cachedata_MPORT_en_pipe_0 = _RAND_1750[0:0];
  _RAND_1751 = {1{`RANDOM}};
  dataArray_36_7_cachedata_MPORT_addr_pipe_0 = _RAND_1751[1:0];
  _RAND_1753 = {1{`RANDOM}};
  dataArray_36_8_cachedata_MPORT_en_pipe_0 = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  dataArray_36_8_cachedata_MPORT_addr_pipe_0 = _RAND_1754[1:0];
  _RAND_1756 = {1{`RANDOM}};
  dataArray_36_9_cachedata_MPORT_en_pipe_0 = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  dataArray_36_9_cachedata_MPORT_addr_pipe_0 = _RAND_1757[1:0];
  _RAND_1759 = {1{`RANDOM}};
  dataArray_36_10_cachedata_MPORT_en_pipe_0 = _RAND_1759[0:0];
  _RAND_1760 = {1{`RANDOM}};
  dataArray_36_10_cachedata_MPORT_addr_pipe_0 = _RAND_1760[1:0];
  _RAND_1762 = {1{`RANDOM}};
  dataArray_36_11_cachedata_MPORT_en_pipe_0 = _RAND_1762[0:0];
  _RAND_1763 = {1{`RANDOM}};
  dataArray_36_11_cachedata_MPORT_addr_pipe_0 = _RAND_1763[1:0];
  _RAND_1765 = {1{`RANDOM}};
  dataArray_36_12_cachedata_MPORT_en_pipe_0 = _RAND_1765[0:0];
  _RAND_1766 = {1{`RANDOM}};
  dataArray_36_12_cachedata_MPORT_addr_pipe_0 = _RAND_1766[1:0];
  _RAND_1768 = {1{`RANDOM}};
  dataArray_36_13_cachedata_MPORT_en_pipe_0 = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  dataArray_36_13_cachedata_MPORT_addr_pipe_0 = _RAND_1769[1:0];
  _RAND_1771 = {1{`RANDOM}};
  dataArray_36_14_cachedata_MPORT_en_pipe_0 = _RAND_1771[0:0];
  _RAND_1772 = {1{`RANDOM}};
  dataArray_36_14_cachedata_MPORT_addr_pipe_0 = _RAND_1772[1:0];
  _RAND_1774 = {1{`RANDOM}};
  dataArray_36_15_cachedata_MPORT_en_pipe_0 = _RAND_1774[0:0];
  _RAND_1775 = {1{`RANDOM}};
  dataArray_36_15_cachedata_MPORT_addr_pipe_0 = _RAND_1775[1:0];
  _RAND_1777 = {1{`RANDOM}};
  dataArray_37_0_cachedata_MPORT_en_pipe_0 = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  dataArray_37_0_cachedata_MPORT_addr_pipe_0 = _RAND_1778[1:0];
  _RAND_1780 = {1{`RANDOM}};
  dataArray_37_1_cachedata_MPORT_en_pipe_0 = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  dataArray_37_1_cachedata_MPORT_addr_pipe_0 = _RAND_1781[1:0];
  _RAND_1783 = {1{`RANDOM}};
  dataArray_37_2_cachedata_MPORT_en_pipe_0 = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  dataArray_37_2_cachedata_MPORT_addr_pipe_0 = _RAND_1784[1:0];
  _RAND_1786 = {1{`RANDOM}};
  dataArray_37_3_cachedata_MPORT_en_pipe_0 = _RAND_1786[0:0];
  _RAND_1787 = {1{`RANDOM}};
  dataArray_37_3_cachedata_MPORT_addr_pipe_0 = _RAND_1787[1:0];
  _RAND_1789 = {1{`RANDOM}};
  dataArray_37_4_cachedata_MPORT_en_pipe_0 = _RAND_1789[0:0];
  _RAND_1790 = {1{`RANDOM}};
  dataArray_37_4_cachedata_MPORT_addr_pipe_0 = _RAND_1790[1:0];
  _RAND_1792 = {1{`RANDOM}};
  dataArray_37_5_cachedata_MPORT_en_pipe_0 = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  dataArray_37_5_cachedata_MPORT_addr_pipe_0 = _RAND_1793[1:0];
  _RAND_1795 = {1{`RANDOM}};
  dataArray_37_6_cachedata_MPORT_en_pipe_0 = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  dataArray_37_6_cachedata_MPORT_addr_pipe_0 = _RAND_1796[1:0];
  _RAND_1798 = {1{`RANDOM}};
  dataArray_37_7_cachedata_MPORT_en_pipe_0 = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  dataArray_37_7_cachedata_MPORT_addr_pipe_0 = _RAND_1799[1:0];
  _RAND_1801 = {1{`RANDOM}};
  dataArray_37_8_cachedata_MPORT_en_pipe_0 = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  dataArray_37_8_cachedata_MPORT_addr_pipe_0 = _RAND_1802[1:0];
  _RAND_1804 = {1{`RANDOM}};
  dataArray_37_9_cachedata_MPORT_en_pipe_0 = _RAND_1804[0:0];
  _RAND_1805 = {1{`RANDOM}};
  dataArray_37_9_cachedata_MPORT_addr_pipe_0 = _RAND_1805[1:0];
  _RAND_1807 = {1{`RANDOM}};
  dataArray_37_10_cachedata_MPORT_en_pipe_0 = _RAND_1807[0:0];
  _RAND_1808 = {1{`RANDOM}};
  dataArray_37_10_cachedata_MPORT_addr_pipe_0 = _RAND_1808[1:0];
  _RAND_1810 = {1{`RANDOM}};
  dataArray_37_11_cachedata_MPORT_en_pipe_0 = _RAND_1810[0:0];
  _RAND_1811 = {1{`RANDOM}};
  dataArray_37_11_cachedata_MPORT_addr_pipe_0 = _RAND_1811[1:0];
  _RAND_1813 = {1{`RANDOM}};
  dataArray_37_12_cachedata_MPORT_en_pipe_0 = _RAND_1813[0:0];
  _RAND_1814 = {1{`RANDOM}};
  dataArray_37_12_cachedata_MPORT_addr_pipe_0 = _RAND_1814[1:0];
  _RAND_1816 = {1{`RANDOM}};
  dataArray_37_13_cachedata_MPORT_en_pipe_0 = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  dataArray_37_13_cachedata_MPORT_addr_pipe_0 = _RAND_1817[1:0];
  _RAND_1819 = {1{`RANDOM}};
  dataArray_37_14_cachedata_MPORT_en_pipe_0 = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  dataArray_37_14_cachedata_MPORT_addr_pipe_0 = _RAND_1820[1:0];
  _RAND_1822 = {1{`RANDOM}};
  dataArray_37_15_cachedata_MPORT_en_pipe_0 = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  dataArray_37_15_cachedata_MPORT_addr_pipe_0 = _RAND_1823[1:0];
  _RAND_1825 = {1{`RANDOM}};
  dataArray_38_0_cachedata_MPORT_en_pipe_0 = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  dataArray_38_0_cachedata_MPORT_addr_pipe_0 = _RAND_1826[1:0];
  _RAND_1828 = {1{`RANDOM}};
  dataArray_38_1_cachedata_MPORT_en_pipe_0 = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  dataArray_38_1_cachedata_MPORT_addr_pipe_0 = _RAND_1829[1:0];
  _RAND_1831 = {1{`RANDOM}};
  dataArray_38_2_cachedata_MPORT_en_pipe_0 = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  dataArray_38_2_cachedata_MPORT_addr_pipe_0 = _RAND_1832[1:0];
  _RAND_1834 = {1{`RANDOM}};
  dataArray_38_3_cachedata_MPORT_en_pipe_0 = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  dataArray_38_3_cachedata_MPORT_addr_pipe_0 = _RAND_1835[1:0];
  _RAND_1837 = {1{`RANDOM}};
  dataArray_38_4_cachedata_MPORT_en_pipe_0 = _RAND_1837[0:0];
  _RAND_1838 = {1{`RANDOM}};
  dataArray_38_4_cachedata_MPORT_addr_pipe_0 = _RAND_1838[1:0];
  _RAND_1840 = {1{`RANDOM}};
  dataArray_38_5_cachedata_MPORT_en_pipe_0 = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  dataArray_38_5_cachedata_MPORT_addr_pipe_0 = _RAND_1841[1:0];
  _RAND_1843 = {1{`RANDOM}};
  dataArray_38_6_cachedata_MPORT_en_pipe_0 = _RAND_1843[0:0];
  _RAND_1844 = {1{`RANDOM}};
  dataArray_38_6_cachedata_MPORT_addr_pipe_0 = _RAND_1844[1:0];
  _RAND_1846 = {1{`RANDOM}};
  dataArray_38_7_cachedata_MPORT_en_pipe_0 = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  dataArray_38_7_cachedata_MPORT_addr_pipe_0 = _RAND_1847[1:0];
  _RAND_1849 = {1{`RANDOM}};
  dataArray_38_8_cachedata_MPORT_en_pipe_0 = _RAND_1849[0:0];
  _RAND_1850 = {1{`RANDOM}};
  dataArray_38_8_cachedata_MPORT_addr_pipe_0 = _RAND_1850[1:0];
  _RAND_1852 = {1{`RANDOM}};
  dataArray_38_9_cachedata_MPORT_en_pipe_0 = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  dataArray_38_9_cachedata_MPORT_addr_pipe_0 = _RAND_1853[1:0];
  _RAND_1855 = {1{`RANDOM}};
  dataArray_38_10_cachedata_MPORT_en_pipe_0 = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  dataArray_38_10_cachedata_MPORT_addr_pipe_0 = _RAND_1856[1:0];
  _RAND_1858 = {1{`RANDOM}};
  dataArray_38_11_cachedata_MPORT_en_pipe_0 = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  dataArray_38_11_cachedata_MPORT_addr_pipe_0 = _RAND_1859[1:0];
  _RAND_1861 = {1{`RANDOM}};
  dataArray_38_12_cachedata_MPORT_en_pipe_0 = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  dataArray_38_12_cachedata_MPORT_addr_pipe_0 = _RAND_1862[1:0];
  _RAND_1864 = {1{`RANDOM}};
  dataArray_38_13_cachedata_MPORT_en_pipe_0 = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  dataArray_38_13_cachedata_MPORT_addr_pipe_0 = _RAND_1865[1:0];
  _RAND_1867 = {1{`RANDOM}};
  dataArray_38_14_cachedata_MPORT_en_pipe_0 = _RAND_1867[0:0];
  _RAND_1868 = {1{`RANDOM}};
  dataArray_38_14_cachedata_MPORT_addr_pipe_0 = _RAND_1868[1:0];
  _RAND_1870 = {1{`RANDOM}};
  dataArray_38_15_cachedata_MPORT_en_pipe_0 = _RAND_1870[0:0];
  _RAND_1871 = {1{`RANDOM}};
  dataArray_38_15_cachedata_MPORT_addr_pipe_0 = _RAND_1871[1:0];
  _RAND_1873 = {1{`RANDOM}};
  dataArray_39_0_cachedata_MPORT_en_pipe_0 = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  dataArray_39_0_cachedata_MPORT_addr_pipe_0 = _RAND_1874[1:0];
  _RAND_1876 = {1{`RANDOM}};
  dataArray_39_1_cachedata_MPORT_en_pipe_0 = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  dataArray_39_1_cachedata_MPORT_addr_pipe_0 = _RAND_1877[1:0];
  _RAND_1879 = {1{`RANDOM}};
  dataArray_39_2_cachedata_MPORT_en_pipe_0 = _RAND_1879[0:0];
  _RAND_1880 = {1{`RANDOM}};
  dataArray_39_2_cachedata_MPORT_addr_pipe_0 = _RAND_1880[1:0];
  _RAND_1882 = {1{`RANDOM}};
  dataArray_39_3_cachedata_MPORT_en_pipe_0 = _RAND_1882[0:0];
  _RAND_1883 = {1{`RANDOM}};
  dataArray_39_3_cachedata_MPORT_addr_pipe_0 = _RAND_1883[1:0];
  _RAND_1885 = {1{`RANDOM}};
  dataArray_39_4_cachedata_MPORT_en_pipe_0 = _RAND_1885[0:0];
  _RAND_1886 = {1{`RANDOM}};
  dataArray_39_4_cachedata_MPORT_addr_pipe_0 = _RAND_1886[1:0];
  _RAND_1888 = {1{`RANDOM}};
  dataArray_39_5_cachedata_MPORT_en_pipe_0 = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  dataArray_39_5_cachedata_MPORT_addr_pipe_0 = _RAND_1889[1:0];
  _RAND_1891 = {1{`RANDOM}};
  dataArray_39_6_cachedata_MPORT_en_pipe_0 = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  dataArray_39_6_cachedata_MPORT_addr_pipe_0 = _RAND_1892[1:0];
  _RAND_1894 = {1{`RANDOM}};
  dataArray_39_7_cachedata_MPORT_en_pipe_0 = _RAND_1894[0:0];
  _RAND_1895 = {1{`RANDOM}};
  dataArray_39_7_cachedata_MPORT_addr_pipe_0 = _RAND_1895[1:0];
  _RAND_1897 = {1{`RANDOM}};
  dataArray_39_8_cachedata_MPORT_en_pipe_0 = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  dataArray_39_8_cachedata_MPORT_addr_pipe_0 = _RAND_1898[1:0];
  _RAND_1900 = {1{`RANDOM}};
  dataArray_39_9_cachedata_MPORT_en_pipe_0 = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  dataArray_39_9_cachedata_MPORT_addr_pipe_0 = _RAND_1901[1:0];
  _RAND_1903 = {1{`RANDOM}};
  dataArray_39_10_cachedata_MPORT_en_pipe_0 = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  dataArray_39_10_cachedata_MPORT_addr_pipe_0 = _RAND_1904[1:0];
  _RAND_1906 = {1{`RANDOM}};
  dataArray_39_11_cachedata_MPORT_en_pipe_0 = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  dataArray_39_11_cachedata_MPORT_addr_pipe_0 = _RAND_1907[1:0];
  _RAND_1909 = {1{`RANDOM}};
  dataArray_39_12_cachedata_MPORT_en_pipe_0 = _RAND_1909[0:0];
  _RAND_1910 = {1{`RANDOM}};
  dataArray_39_12_cachedata_MPORT_addr_pipe_0 = _RAND_1910[1:0];
  _RAND_1912 = {1{`RANDOM}};
  dataArray_39_13_cachedata_MPORT_en_pipe_0 = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  dataArray_39_13_cachedata_MPORT_addr_pipe_0 = _RAND_1913[1:0];
  _RAND_1915 = {1{`RANDOM}};
  dataArray_39_14_cachedata_MPORT_en_pipe_0 = _RAND_1915[0:0];
  _RAND_1916 = {1{`RANDOM}};
  dataArray_39_14_cachedata_MPORT_addr_pipe_0 = _RAND_1916[1:0];
  _RAND_1918 = {1{`RANDOM}};
  dataArray_39_15_cachedata_MPORT_en_pipe_0 = _RAND_1918[0:0];
  _RAND_1919 = {1{`RANDOM}};
  dataArray_39_15_cachedata_MPORT_addr_pipe_0 = _RAND_1919[1:0];
  _RAND_1921 = {1{`RANDOM}};
  dataArray_40_0_cachedata_MPORT_en_pipe_0 = _RAND_1921[0:0];
  _RAND_1922 = {1{`RANDOM}};
  dataArray_40_0_cachedata_MPORT_addr_pipe_0 = _RAND_1922[1:0];
  _RAND_1924 = {1{`RANDOM}};
  dataArray_40_1_cachedata_MPORT_en_pipe_0 = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  dataArray_40_1_cachedata_MPORT_addr_pipe_0 = _RAND_1925[1:0];
  _RAND_1927 = {1{`RANDOM}};
  dataArray_40_2_cachedata_MPORT_en_pipe_0 = _RAND_1927[0:0];
  _RAND_1928 = {1{`RANDOM}};
  dataArray_40_2_cachedata_MPORT_addr_pipe_0 = _RAND_1928[1:0];
  _RAND_1930 = {1{`RANDOM}};
  dataArray_40_3_cachedata_MPORT_en_pipe_0 = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  dataArray_40_3_cachedata_MPORT_addr_pipe_0 = _RAND_1931[1:0];
  _RAND_1933 = {1{`RANDOM}};
  dataArray_40_4_cachedata_MPORT_en_pipe_0 = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  dataArray_40_4_cachedata_MPORT_addr_pipe_0 = _RAND_1934[1:0];
  _RAND_1936 = {1{`RANDOM}};
  dataArray_40_5_cachedata_MPORT_en_pipe_0 = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  dataArray_40_5_cachedata_MPORT_addr_pipe_0 = _RAND_1937[1:0];
  _RAND_1939 = {1{`RANDOM}};
  dataArray_40_6_cachedata_MPORT_en_pipe_0 = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  dataArray_40_6_cachedata_MPORT_addr_pipe_0 = _RAND_1940[1:0];
  _RAND_1942 = {1{`RANDOM}};
  dataArray_40_7_cachedata_MPORT_en_pipe_0 = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  dataArray_40_7_cachedata_MPORT_addr_pipe_0 = _RAND_1943[1:0];
  _RAND_1945 = {1{`RANDOM}};
  dataArray_40_8_cachedata_MPORT_en_pipe_0 = _RAND_1945[0:0];
  _RAND_1946 = {1{`RANDOM}};
  dataArray_40_8_cachedata_MPORT_addr_pipe_0 = _RAND_1946[1:0];
  _RAND_1948 = {1{`RANDOM}};
  dataArray_40_9_cachedata_MPORT_en_pipe_0 = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  dataArray_40_9_cachedata_MPORT_addr_pipe_0 = _RAND_1949[1:0];
  _RAND_1951 = {1{`RANDOM}};
  dataArray_40_10_cachedata_MPORT_en_pipe_0 = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  dataArray_40_10_cachedata_MPORT_addr_pipe_0 = _RAND_1952[1:0];
  _RAND_1954 = {1{`RANDOM}};
  dataArray_40_11_cachedata_MPORT_en_pipe_0 = _RAND_1954[0:0];
  _RAND_1955 = {1{`RANDOM}};
  dataArray_40_11_cachedata_MPORT_addr_pipe_0 = _RAND_1955[1:0];
  _RAND_1957 = {1{`RANDOM}};
  dataArray_40_12_cachedata_MPORT_en_pipe_0 = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  dataArray_40_12_cachedata_MPORT_addr_pipe_0 = _RAND_1958[1:0];
  _RAND_1960 = {1{`RANDOM}};
  dataArray_40_13_cachedata_MPORT_en_pipe_0 = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  dataArray_40_13_cachedata_MPORT_addr_pipe_0 = _RAND_1961[1:0];
  _RAND_1963 = {1{`RANDOM}};
  dataArray_40_14_cachedata_MPORT_en_pipe_0 = _RAND_1963[0:0];
  _RAND_1964 = {1{`RANDOM}};
  dataArray_40_14_cachedata_MPORT_addr_pipe_0 = _RAND_1964[1:0];
  _RAND_1966 = {1{`RANDOM}};
  dataArray_40_15_cachedata_MPORT_en_pipe_0 = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  dataArray_40_15_cachedata_MPORT_addr_pipe_0 = _RAND_1967[1:0];
  _RAND_1969 = {1{`RANDOM}};
  dataArray_41_0_cachedata_MPORT_en_pipe_0 = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  dataArray_41_0_cachedata_MPORT_addr_pipe_0 = _RAND_1970[1:0];
  _RAND_1972 = {1{`RANDOM}};
  dataArray_41_1_cachedata_MPORT_en_pipe_0 = _RAND_1972[0:0];
  _RAND_1973 = {1{`RANDOM}};
  dataArray_41_1_cachedata_MPORT_addr_pipe_0 = _RAND_1973[1:0];
  _RAND_1975 = {1{`RANDOM}};
  dataArray_41_2_cachedata_MPORT_en_pipe_0 = _RAND_1975[0:0];
  _RAND_1976 = {1{`RANDOM}};
  dataArray_41_2_cachedata_MPORT_addr_pipe_0 = _RAND_1976[1:0];
  _RAND_1978 = {1{`RANDOM}};
  dataArray_41_3_cachedata_MPORT_en_pipe_0 = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  dataArray_41_3_cachedata_MPORT_addr_pipe_0 = _RAND_1979[1:0];
  _RAND_1981 = {1{`RANDOM}};
  dataArray_41_4_cachedata_MPORT_en_pipe_0 = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  dataArray_41_4_cachedata_MPORT_addr_pipe_0 = _RAND_1982[1:0];
  _RAND_1984 = {1{`RANDOM}};
  dataArray_41_5_cachedata_MPORT_en_pipe_0 = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  dataArray_41_5_cachedata_MPORT_addr_pipe_0 = _RAND_1985[1:0];
  _RAND_1987 = {1{`RANDOM}};
  dataArray_41_6_cachedata_MPORT_en_pipe_0 = _RAND_1987[0:0];
  _RAND_1988 = {1{`RANDOM}};
  dataArray_41_6_cachedata_MPORT_addr_pipe_0 = _RAND_1988[1:0];
  _RAND_1990 = {1{`RANDOM}};
  dataArray_41_7_cachedata_MPORT_en_pipe_0 = _RAND_1990[0:0];
  _RAND_1991 = {1{`RANDOM}};
  dataArray_41_7_cachedata_MPORT_addr_pipe_0 = _RAND_1991[1:0];
  _RAND_1993 = {1{`RANDOM}};
  dataArray_41_8_cachedata_MPORT_en_pipe_0 = _RAND_1993[0:0];
  _RAND_1994 = {1{`RANDOM}};
  dataArray_41_8_cachedata_MPORT_addr_pipe_0 = _RAND_1994[1:0];
  _RAND_1996 = {1{`RANDOM}};
  dataArray_41_9_cachedata_MPORT_en_pipe_0 = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  dataArray_41_9_cachedata_MPORT_addr_pipe_0 = _RAND_1997[1:0];
  _RAND_1999 = {1{`RANDOM}};
  dataArray_41_10_cachedata_MPORT_en_pipe_0 = _RAND_1999[0:0];
  _RAND_2000 = {1{`RANDOM}};
  dataArray_41_10_cachedata_MPORT_addr_pipe_0 = _RAND_2000[1:0];
  _RAND_2002 = {1{`RANDOM}};
  dataArray_41_11_cachedata_MPORT_en_pipe_0 = _RAND_2002[0:0];
  _RAND_2003 = {1{`RANDOM}};
  dataArray_41_11_cachedata_MPORT_addr_pipe_0 = _RAND_2003[1:0];
  _RAND_2005 = {1{`RANDOM}};
  dataArray_41_12_cachedata_MPORT_en_pipe_0 = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  dataArray_41_12_cachedata_MPORT_addr_pipe_0 = _RAND_2006[1:0];
  _RAND_2008 = {1{`RANDOM}};
  dataArray_41_13_cachedata_MPORT_en_pipe_0 = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  dataArray_41_13_cachedata_MPORT_addr_pipe_0 = _RAND_2009[1:0];
  _RAND_2011 = {1{`RANDOM}};
  dataArray_41_14_cachedata_MPORT_en_pipe_0 = _RAND_2011[0:0];
  _RAND_2012 = {1{`RANDOM}};
  dataArray_41_14_cachedata_MPORT_addr_pipe_0 = _RAND_2012[1:0];
  _RAND_2014 = {1{`RANDOM}};
  dataArray_41_15_cachedata_MPORT_en_pipe_0 = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  dataArray_41_15_cachedata_MPORT_addr_pipe_0 = _RAND_2015[1:0];
  _RAND_2017 = {1{`RANDOM}};
  dataArray_42_0_cachedata_MPORT_en_pipe_0 = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  dataArray_42_0_cachedata_MPORT_addr_pipe_0 = _RAND_2018[1:0];
  _RAND_2020 = {1{`RANDOM}};
  dataArray_42_1_cachedata_MPORT_en_pipe_0 = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  dataArray_42_1_cachedata_MPORT_addr_pipe_0 = _RAND_2021[1:0];
  _RAND_2023 = {1{`RANDOM}};
  dataArray_42_2_cachedata_MPORT_en_pipe_0 = _RAND_2023[0:0];
  _RAND_2024 = {1{`RANDOM}};
  dataArray_42_2_cachedata_MPORT_addr_pipe_0 = _RAND_2024[1:0];
  _RAND_2026 = {1{`RANDOM}};
  dataArray_42_3_cachedata_MPORT_en_pipe_0 = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  dataArray_42_3_cachedata_MPORT_addr_pipe_0 = _RAND_2027[1:0];
  _RAND_2029 = {1{`RANDOM}};
  dataArray_42_4_cachedata_MPORT_en_pipe_0 = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  dataArray_42_4_cachedata_MPORT_addr_pipe_0 = _RAND_2030[1:0];
  _RAND_2032 = {1{`RANDOM}};
  dataArray_42_5_cachedata_MPORT_en_pipe_0 = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  dataArray_42_5_cachedata_MPORT_addr_pipe_0 = _RAND_2033[1:0];
  _RAND_2035 = {1{`RANDOM}};
  dataArray_42_6_cachedata_MPORT_en_pipe_0 = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  dataArray_42_6_cachedata_MPORT_addr_pipe_0 = _RAND_2036[1:0];
  _RAND_2038 = {1{`RANDOM}};
  dataArray_42_7_cachedata_MPORT_en_pipe_0 = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  dataArray_42_7_cachedata_MPORT_addr_pipe_0 = _RAND_2039[1:0];
  _RAND_2041 = {1{`RANDOM}};
  dataArray_42_8_cachedata_MPORT_en_pipe_0 = _RAND_2041[0:0];
  _RAND_2042 = {1{`RANDOM}};
  dataArray_42_8_cachedata_MPORT_addr_pipe_0 = _RAND_2042[1:0];
  _RAND_2044 = {1{`RANDOM}};
  dataArray_42_9_cachedata_MPORT_en_pipe_0 = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  dataArray_42_9_cachedata_MPORT_addr_pipe_0 = _RAND_2045[1:0];
  _RAND_2047 = {1{`RANDOM}};
  dataArray_42_10_cachedata_MPORT_en_pipe_0 = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  dataArray_42_10_cachedata_MPORT_addr_pipe_0 = _RAND_2048[1:0];
  _RAND_2050 = {1{`RANDOM}};
  dataArray_42_11_cachedata_MPORT_en_pipe_0 = _RAND_2050[0:0];
  _RAND_2051 = {1{`RANDOM}};
  dataArray_42_11_cachedata_MPORT_addr_pipe_0 = _RAND_2051[1:0];
  _RAND_2053 = {1{`RANDOM}};
  dataArray_42_12_cachedata_MPORT_en_pipe_0 = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  dataArray_42_12_cachedata_MPORT_addr_pipe_0 = _RAND_2054[1:0];
  _RAND_2056 = {1{`RANDOM}};
  dataArray_42_13_cachedata_MPORT_en_pipe_0 = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  dataArray_42_13_cachedata_MPORT_addr_pipe_0 = _RAND_2057[1:0];
  _RAND_2059 = {1{`RANDOM}};
  dataArray_42_14_cachedata_MPORT_en_pipe_0 = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  dataArray_42_14_cachedata_MPORT_addr_pipe_0 = _RAND_2060[1:0];
  _RAND_2062 = {1{`RANDOM}};
  dataArray_42_15_cachedata_MPORT_en_pipe_0 = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  dataArray_42_15_cachedata_MPORT_addr_pipe_0 = _RAND_2063[1:0];
  _RAND_2065 = {1{`RANDOM}};
  dataArray_43_0_cachedata_MPORT_en_pipe_0 = _RAND_2065[0:0];
  _RAND_2066 = {1{`RANDOM}};
  dataArray_43_0_cachedata_MPORT_addr_pipe_0 = _RAND_2066[1:0];
  _RAND_2068 = {1{`RANDOM}};
  dataArray_43_1_cachedata_MPORT_en_pipe_0 = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  dataArray_43_1_cachedata_MPORT_addr_pipe_0 = _RAND_2069[1:0];
  _RAND_2071 = {1{`RANDOM}};
  dataArray_43_2_cachedata_MPORT_en_pipe_0 = _RAND_2071[0:0];
  _RAND_2072 = {1{`RANDOM}};
  dataArray_43_2_cachedata_MPORT_addr_pipe_0 = _RAND_2072[1:0];
  _RAND_2074 = {1{`RANDOM}};
  dataArray_43_3_cachedata_MPORT_en_pipe_0 = _RAND_2074[0:0];
  _RAND_2075 = {1{`RANDOM}};
  dataArray_43_3_cachedata_MPORT_addr_pipe_0 = _RAND_2075[1:0];
  _RAND_2077 = {1{`RANDOM}};
  dataArray_43_4_cachedata_MPORT_en_pipe_0 = _RAND_2077[0:0];
  _RAND_2078 = {1{`RANDOM}};
  dataArray_43_4_cachedata_MPORT_addr_pipe_0 = _RAND_2078[1:0];
  _RAND_2080 = {1{`RANDOM}};
  dataArray_43_5_cachedata_MPORT_en_pipe_0 = _RAND_2080[0:0];
  _RAND_2081 = {1{`RANDOM}};
  dataArray_43_5_cachedata_MPORT_addr_pipe_0 = _RAND_2081[1:0];
  _RAND_2083 = {1{`RANDOM}};
  dataArray_43_6_cachedata_MPORT_en_pipe_0 = _RAND_2083[0:0];
  _RAND_2084 = {1{`RANDOM}};
  dataArray_43_6_cachedata_MPORT_addr_pipe_0 = _RAND_2084[1:0];
  _RAND_2086 = {1{`RANDOM}};
  dataArray_43_7_cachedata_MPORT_en_pipe_0 = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  dataArray_43_7_cachedata_MPORT_addr_pipe_0 = _RAND_2087[1:0];
  _RAND_2089 = {1{`RANDOM}};
  dataArray_43_8_cachedata_MPORT_en_pipe_0 = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  dataArray_43_8_cachedata_MPORT_addr_pipe_0 = _RAND_2090[1:0];
  _RAND_2092 = {1{`RANDOM}};
  dataArray_43_9_cachedata_MPORT_en_pipe_0 = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  dataArray_43_9_cachedata_MPORT_addr_pipe_0 = _RAND_2093[1:0];
  _RAND_2095 = {1{`RANDOM}};
  dataArray_43_10_cachedata_MPORT_en_pipe_0 = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  dataArray_43_10_cachedata_MPORT_addr_pipe_0 = _RAND_2096[1:0];
  _RAND_2098 = {1{`RANDOM}};
  dataArray_43_11_cachedata_MPORT_en_pipe_0 = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  dataArray_43_11_cachedata_MPORT_addr_pipe_0 = _RAND_2099[1:0];
  _RAND_2101 = {1{`RANDOM}};
  dataArray_43_12_cachedata_MPORT_en_pipe_0 = _RAND_2101[0:0];
  _RAND_2102 = {1{`RANDOM}};
  dataArray_43_12_cachedata_MPORT_addr_pipe_0 = _RAND_2102[1:0];
  _RAND_2104 = {1{`RANDOM}};
  dataArray_43_13_cachedata_MPORT_en_pipe_0 = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  dataArray_43_13_cachedata_MPORT_addr_pipe_0 = _RAND_2105[1:0];
  _RAND_2107 = {1{`RANDOM}};
  dataArray_43_14_cachedata_MPORT_en_pipe_0 = _RAND_2107[0:0];
  _RAND_2108 = {1{`RANDOM}};
  dataArray_43_14_cachedata_MPORT_addr_pipe_0 = _RAND_2108[1:0];
  _RAND_2110 = {1{`RANDOM}};
  dataArray_43_15_cachedata_MPORT_en_pipe_0 = _RAND_2110[0:0];
  _RAND_2111 = {1{`RANDOM}};
  dataArray_43_15_cachedata_MPORT_addr_pipe_0 = _RAND_2111[1:0];
  _RAND_2113 = {1{`RANDOM}};
  dataArray_44_0_cachedata_MPORT_en_pipe_0 = _RAND_2113[0:0];
  _RAND_2114 = {1{`RANDOM}};
  dataArray_44_0_cachedata_MPORT_addr_pipe_0 = _RAND_2114[1:0];
  _RAND_2116 = {1{`RANDOM}};
  dataArray_44_1_cachedata_MPORT_en_pipe_0 = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  dataArray_44_1_cachedata_MPORT_addr_pipe_0 = _RAND_2117[1:0];
  _RAND_2119 = {1{`RANDOM}};
  dataArray_44_2_cachedata_MPORT_en_pipe_0 = _RAND_2119[0:0];
  _RAND_2120 = {1{`RANDOM}};
  dataArray_44_2_cachedata_MPORT_addr_pipe_0 = _RAND_2120[1:0];
  _RAND_2122 = {1{`RANDOM}};
  dataArray_44_3_cachedata_MPORT_en_pipe_0 = _RAND_2122[0:0];
  _RAND_2123 = {1{`RANDOM}};
  dataArray_44_3_cachedata_MPORT_addr_pipe_0 = _RAND_2123[1:0];
  _RAND_2125 = {1{`RANDOM}};
  dataArray_44_4_cachedata_MPORT_en_pipe_0 = _RAND_2125[0:0];
  _RAND_2126 = {1{`RANDOM}};
  dataArray_44_4_cachedata_MPORT_addr_pipe_0 = _RAND_2126[1:0];
  _RAND_2128 = {1{`RANDOM}};
  dataArray_44_5_cachedata_MPORT_en_pipe_0 = _RAND_2128[0:0];
  _RAND_2129 = {1{`RANDOM}};
  dataArray_44_5_cachedata_MPORT_addr_pipe_0 = _RAND_2129[1:0];
  _RAND_2131 = {1{`RANDOM}};
  dataArray_44_6_cachedata_MPORT_en_pipe_0 = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  dataArray_44_6_cachedata_MPORT_addr_pipe_0 = _RAND_2132[1:0];
  _RAND_2134 = {1{`RANDOM}};
  dataArray_44_7_cachedata_MPORT_en_pipe_0 = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  dataArray_44_7_cachedata_MPORT_addr_pipe_0 = _RAND_2135[1:0];
  _RAND_2137 = {1{`RANDOM}};
  dataArray_44_8_cachedata_MPORT_en_pipe_0 = _RAND_2137[0:0];
  _RAND_2138 = {1{`RANDOM}};
  dataArray_44_8_cachedata_MPORT_addr_pipe_0 = _RAND_2138[1:0];
  _RAND_2140 = {1{`RANDOM}};
  dataArray_44_9_cachedata_MPORT_en_pipe_0 = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  dataArray_44_9_cachedata_MPORT_addr_pipe_0 = _RAND_2141[1:0];
  _RAND_2143 = {1{`RANDOM}};
  dataArray_44_10_cachedata_MPORT_en_pipe_0 = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  dataArray_44_10_cachedata_MPORT_addr_pipe_0 = _RAND_2144[1:0];
  _RAND_2146 = {1{`RANDOM}};
  dataArray_44_11_cachedata_MPORT_en_pipe_0 = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  dataArray_44_11_cachedata_MPORT_addr_pipe_0 = _RAND_2147[1:0];
  _RAND_2149 = {1{`RANDOM}};
  dataArray_44_12_cachedata_MPORT_en_pipe_0 = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  dataArray_44_12_cachedata_MPORT_addr_pipe_0 = _RAND_2150[1:0];
  _RAND_2152 = {1{`RANDOM}};
  dataArray_44_13_cachedata_MPORT_en_pipe_0 = _RAND_2152[0:0];
  _RAND_2153 = {1{`RANDOM}};
  dataArray_44_13_cachedata_MPORT_addr_pipe_0 = _RAND_2153[1:0];
  _RAND_2155 = {1{`RANDOM}};
  dataArray_44_14_cachedata_MPORT_en_pipe_0 = _RAND_2155[0:0];
  _RAND_2156 = {1{`RANDOM}};
  dataArray_44_14_cachedata_MPORT_addr_pipe_0 = _RAND_2156[1:0];
  _RAND_2158 = {1{`RANDOM}};
  dataArray_44_15_cachedata_MPORT_en_pipe_0 = _RAND_2158[0:0];
  _RAND_2159 = {1{`RANDOM}};
  dataArray_44_15_cachedata_MPORT_addr_pipe_0 = _RAND_2159[1:0];
  _RAND_2161 = {1{`RANDOM}};
  dataArray_45_0_cachedata_MPORT_en_pipe_0 = _RAND_2161[0:0];
  _RAND_2162 = {1{`RANDOM}};
  dataArray_45_0_cachedata_MPORT_addr_pipe_0 = _RAND_2162[1:0];
  _RAND_2164 = {1{`RANDOM}};
  dataArray_45_1_cachedata_MPORT_en_pipe_0 = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  dataArray_45_1_cachedata_MPORT_addr_pipe_0 = _RAND_2165[1:0];
  _RAND_2167 = {1{`RANDOM}};
  dataArray_45_2_cachedata_MPORT_en_pipe_0 = _RAND_2167[0:0];
  _RAND_2168 = {1{`RANDOM}};
  dataArray_45_2_cachedata_MPORT_addr_pipe_0 = _RAND_2168[1:0];
  _RAND_2170 = {1{`RANDOM}};
  dataArray_45_3_cachedata_MPORT_en_pipe_0 = _RAND_2170[0:0];
  _RAND_2171 = {1{`RANDOM}};
  dataArray_45_3_cachedata_MPORT_addr_pipe_0 = _RAND_2171[1:0];
  _RAND_2173 = {1{`RANDOM}};
  dataArray_45_4_cachedata_MPORT_en_pipe_0 = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  dataArray_45_4_cachedata_MPORT_addr_pipe_0 = _RAND_2174[1:0];
  _RAND_2176 = {1{`RANDOM}};
  dataArray_45_5_cachedata_MPORT_en_pipe_0 = _RAND_2176[0:0];
  _RAND_2177 = {1{`RANDOM}};
  dataArray_45_5_cachedata_MPORT_addr_pipe_0 = _RAND_2177[1:0];
  _RAND_2179 = {1{`RANDOM}};
  dataArray_45_6_cachedata_MPORT_en_pipe_0 = _RAND_2179[0:0];
  _RAND_2180 = {1{`RANDOM}};
  dataArray_45_6_cachedata_MPORT_addr_pipe_0 = _RAND_2180[1:0];
  _RAND_2182 = {1{`RANDOM}};
  dataArray_45_7_cachedata_MPORT_en_pipe_0 = _RAND_2182[0:0];
  _RAND_2183 = {1{`RANDOM}};
  dataArray_45_7_cachedata_MPORT_addr_pipe_0 = _RAND_2183[1:0];
  _RAND_2185 = {1{`RANDOM}};
  dataArray_45_8_cachedata_MPORT_en_pipe_0 = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  dataArray_45_8_cachedata_MPORT_addr_pipe_0 = _RAND_2186[1:0];
  _RAND_2188 = {1{`RANDOM}};
  dataArray_45_9_cachedata_MPORT_en_pipe_0 = _RAND_2188[0:0];
  _RAND_2189 = {1{`RANDOM}};
  dataArray_45_9_cachedata_MPORT_addr_pipe_0 = _RAND_2189[1:0];
  _RAND_2191 = {1{`RANDOM}};
  dataArray_45_10_cachedata_MPORT_en_pipe_0 = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  dataArray_45_10_cachedata_MPORT_addr_pipe_0 = _RAND_2192[1:0];
  _RAND_2194 = {1{`RANDOM}};
  dataArray_45_11_cachedata_MPORT_en_pipe_0 = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  dataArray_45_11_cachedata_MPORT_addr_pipe_0 = _RAND_2195[1:0];
  _RAND_2197 = {1{`RANDOM}};
  dataArray_45_12_cachedata_MPORT_en_pipe_0 = _RAND_2197[0:0];
  _RAND_2198 = {1{`RANDOM}};
  dataArray_45_12_cachedata_MPORT_addr_pipe_0 = _RAND_2198[1:0];
  _RAND_2200 = {1{`RANDOM}};
  dataArray_45_13_cachedata_MPORT_en_pipe_0 = _RAND_2200[0:0];
  _RAND_2201 = {1{`RANDOM}};
  dataArray_45_13_cachedata_MPORT_addr_pipe_0 = _RAND_2201[1:0];
  _RAND_2203 = {1{`RANDOM}};
  dataArray_45_14_cachedata_MPORT_en_pipe_0 = _RAND_2203[0:0];
  _RAND_2204 = {1{`RANDOM}};
  dataArray_45_14_cachedata_MPORT_addr_pipe_0 = _RAND_2204[1:0];
  _RAND_2206 = {1{`RANDOM}};
  dataArray_45_15_cachedata_MPORT_en_pipe_0 = _RAND_2206[0:0];
  _RAND_2207 = {1{`RANDOM}};
  dataArray_45_15_cachedata_MPORT_addr_pipe_0 = _RAND_2207[1:0];
  _RAND_2209 = {1{`RANDOM}};
  dataArray_46_0_cachedata_MPORT_en_pipe_0 = _RAND_2209[0:0];
  _RAND_2210 = {1{`RANDOM}};
  dataArray_46_0_cachedata_MPORT_addr_pipe_0 = _RAND_2210[1:0];
  _RAND_2212 = {1{`RANDOM}};
  dataArray_46_1_cachedata_MPORT_en_pipe_0 = _RAND_2212[0:0];
  _RAND_2213 = {1{`RANDOM}};
  dataArray_46_1_cachedata_MPORT_addr_pipe_0 = _RAND_2213[1:0];
  _RAND_2215 = {1{`RANDOM}};
  dataArray_46_2_cachedata_MPORT_en_pipe_0 = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  dataArray_46_2_cachedata_MPORT_addr_pipe_0 = _RAND_2216[1:0];
  _RAND_2218 = {1{`RANDOM}};
  dataArray_46_3_cachedata_MPORT_en_pipe_0 = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  dataArray_46_3_cachedata_MPORT_addr_pipe_0 = _RAND_2219[1:0];
  _RAND_2221 = {1{`RANDOM}};
  dataArray_46_4_cachedata_MPORT_en_pipe_0 = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  dataArray_46_4_cachedata_MPORT_addr_pipe_0 = _RAND_2222[1:0];
  _RAND_2224 = {1{`RANDOM}};
  dataArray_46_5_cachedata_MPORT_en_pipe_0 = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  dataArray_46_5_cachedata_MPORT_addr_pipe_0 = _RAND_2225[1:0];
  _RAND_2227 = {1{`RANDOM}};
  dataArray_46_6_cachedata_MPORT_en_pipe_0 = _RAND_2227[0:0];
  _RAND_2228 = {1{`RANDOM}};
  dataArray_46_6_cachedata_MPORT_addr_pipe_0 = _RAND_2228[1:0];
  _RAND_2230 = {1{`RANDOM}};
  dataArray_46_7_cachedata_MPORT_en_pipe_0 = _RAND_2230[0:0];
  _RAND_2231 = {1{`RANDOM}};
  dataArray_46_7_cachedata_MPORT_addr_pipe_0 = _RAND_2231[1:0];
  _RAND_2233 = {1{`RANDOM}};
  dataArray_46_8_cachedata_MPORT_en_pipe_0 = _RAND_2233[0:0];
  _RAND_2234 = {1{`RANDOM}};
  dataArray_46_8_cachedata_MPORT_addr_pipe_0 = _RAND_2234[1:0];
  _RAND_2236 = {1{`RANDOM}};
  dataArray_46_9_cachedata_MPORT_en_pipe_0 = _RAND_2236[0:0];
  _RAND_2237 = {1{`RANDOM}};
  dataArray_46_9_cachedata_MPORT_addr_pipe_0 = _RAND_2237[1:0];
  _RAND_2239 = {1{`RANDOM}};
  dataArray_46_10_cachedata_MPORT_en_pipe_0 = _RAND_2239[0:0];
  _RAND_2240 = {1{`RANDOM}};
  dataArray_46_10_cachedata_MPORT_addr_pipe_0 = _RAND_2240[1:0];
  _RAND_2242 = {1{`RANDOM}};
  dataArray_46_11_cachedata_MPORT_en_pipe_0 = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  dataArray_46_11_cachedata_MPORT_addr_pipe_0 = _RAND_2243[1:0];
  _RAND_2245 = {1{`RANDOM}};
  dataArray_46_12_cachedata_MPORT_en_pipe_0 = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  dataArray_46_12_cachedata_MPORT_addr_pipe_0 = _RAND_2246[1:0];
  _RAND_2248 = {1{`RANDOM}};
  dataArray_46_13_cachedata_MPORT_en_pipe_0 = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  dataArray_46_13_cachedata_MPORT_addr_pipe_0 = _RAND_2249[1:0];
  _RAND_2251 = {1{`RANDOM}};
  dataArray_46_14_cachedata_MPORT_en_pipe_0 = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  dataArray_46_14_cachedata_MPORT_addr_pipe_0 = _RAND_2252[1:0];
  _RAND_2254 = {1{`RANDOM}};
  dataArray_46_15_cachedata_MPORT_en_pipe_0 = _RAND_2254[0:0];
  _RAND_2255 = {1{`RANDOM}};
  dataArray_46_15_cachedata_MPORT_addr_pipe_0 = _RAND_2255[1:0];
  _RAND_2257 = {1{`RANDOM}};
  dataArray_47_0_cachedata_MPORT_en_pipe_0 = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  dataArray_47_0_cachedata_MPORT_addr_pipe_0 = _RAND_2258[1:0];
  _RAND_2260 = {1{`RANDOM}};
  dataArray_47_1_cachedata_MPORT_en_pipe_0 = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  dataArray_47_1_cachedata_MPORT_addr_pipe_0 = _RAND_2261[1:0];
  _RAND_2263 = {1{`RANDOM}};
  dataArray_47_2_cachedata_MPORT_en_pipe_0 = _RAND_2263[0:0];
  _RAND_2264 = {1{`RANDOM}};
  dataArray_47_2_cachedata_MPORT_addr_pipe_0 = _RAND_2264[1:0];
  _RAND_2266 = {1{`RANDOM}};
  dataArray_47_3_cachedata_MPORT_en_pipe_0 = _RAND_2266[0:0];
  _RAND_2267 = {1{`RANDOM}};
  dataArray_47_3_cachedata_MPORT_addr_pipe_0 = _RAND_2267[1:0];
  _RAND_2269 = {1{`RANDOM}};
  dataArray_47_4_cachedata_MPORT_en_pipe_0 = _RAND_2269[0:0];
  _RAND_2270 = {1{`RANDOM}};
  dataArray_47_4_cachedata_MPORT_addr_pipe_0 = _RAND_2270[1:0];
  _RAND_2272 = {1{`RANDOM}};
  dataArray_47_5_cachedata_MPORT_en_pipe_0 = _RAND_2272[0:0];
  _RAND_2273 = {1{`RANDOM}};
  dataArray_47_5_cachedata_MPORT_addr_pipe_0 = _RAND_2273[1:0];
  _RAND_2275 = {1{`RANDOM}};
  dataArray_47_6_cachedata_MPORT_en_pipe_0 = _RAND_2275[0:0];
  _RAND_2276 = {1{`RANDOM}};
  dataArray_47_6_cachedata_MPORT_addr_pipe_0 = _RAND_2276[1:0];
  _RAND_2278 = {1{`RANDOM}};
  dataArray_47_7_cachedata_MPORT_en_pipe_0 = _RAND_2278[0:0];
  _RAND_2279 = {1{`RANDOM}};
  dataArray_47_7_cachedata_MPORT_addr_pipe_0 = _RAND_2279[1:0];
  _RAND_2281 = {1{`RANDOM}};
  dataArray_47_8_cachedata_MPORT_en_pipe_0 = _RAND_2281[0:0];
  _RAND_2282 = {1{`RANDOM}};
  dataArray_47_8_cachedata_MPORT_addr_pipe_0 = _RAND_2282[1:0];
  _RAND_2284 = {1{`RANDOM}};
  dataArray_47_9_cachedata_MPORT_en_pipe_0 = _RAND_2284[0:0];
  _RAND_2285 = {1{`RANDOM}};
  dataArray_47_9_cachedata_MPORT_addr_pipe_0 = _RAND_2285[1:0];
  _RAND_2287 = {1{`RANDOM}};
  dataArray_47_10_cachedata_MPORT_en_pipe_0 = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  dataArray_47_10_cachedata_MPORT_addr_pipe_0 = _RAND_2288[1:0];
  _RAND_2290 = {1{`RANDOM}};
  dataArray_47_11_cachedata_MPORT_en_pipe_0 = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  dataArray_47_11_cachedata_MPORT_addr_pipe_0 = _RAND_2291[1:0];
  _RAND_2293 = {1{`RANDOM}};
  dataArray_47_12_cachedata_MPORT_en_pipe_0 = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  dataArray_47_12_cachedata_MPORT_addr_pipe_0 = _RAND_2294[1:0];
  _RAND_2296 = {1{`RANDOM}};
  dataArray_47_13_cachedata_MPORT_en_pipe_0 = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  dataArray_47_13_cachedata_MPORT_addr_pipe_0 = _RAND_2297[1:0];
  _RAND_2299 = {1{`RANDOM}};
  dataArray_47_14_cachedata_MPORT_en_pipe_0 = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  dataArray_47_14_cachedata_MPORT_addr_pipe_0 = _RAND_2300[1:0];
  _RAND_2302 = {1{`RANDOM}};
  dataArray_47_15_cachedata_MPORT_en_pipe_0 = _RAND_2302[0:0];
  _RAND_2303 = {1{`RANDOM}};
  dataArray_47_15_cachedata_MPORT_addr_pipe_0 = _RAND_2303[1:0];
  _RAND_2305 = {1{`RANDOM}};
  dataArray_48_0_cachedata_MPORT_en_pipe_0 = _RAND_2305[0:0];
  _RAND_2306 = {1{`RANDOM}};
  dataArray_48_0_cachedata_MPORT_addr_pipe_0 = _RAND_2306[1:0];
  _RAND_2308 = {1{`RANDOM}};
  dataArray_48_1_cachedata_MPORT_en_pipe_0 = _RAND_2308[0:0];
  _RAND_2309 = {1{`RANDOM}};
  dataArray_48_1_cachedata_MPORT_addr_pipe_0 = _RAND_2309[1:0];
  _RAND_2311 = {1{`RANDOM}};
  dataArray_48_2_cachedata_MPORT_en_pipe_0 = _RAND_2311[0:0];
  _RAND_2312 = {1{`RANDOM}};
  dataArray_48_2_cachedata_MPORT_addr_pipe_0 = _RAND_2312[1:0];
  _RAND_2314 = {1{`RANDOM}};
  dataArray_48_3_cachedata_MPORT_en_pipe_0 = _RAND_2314[0:0];
  _RAND_2315 = {1{`RANDOM}};
  dataArray_48_3_cachedata_MPORT_addr_pipe_0 = _RAND_2315[1:0];
  _RAND_2317 = {1{`RANDOM}};
  dataArray_48_4_cachedata_MPORT_en_pipe_0 = _RAND_2317[0:0];
  _RAND_2318 = {1{`RANDOM}};
  dataArray_48_4_cachedata_MPORT_addr_pipe_0 = _RAND_2318[1:0];
  _RAND_2320 = {1{`RANDOM}};
  dataArray_48_5_cachedata_MPORT_en_pipe_0 = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  dataArray_48_5_cachedata_MPORT_addr_pipe_0 = _RAND_2321[1:0];
  _RAND_2323 = {1{`RANDOM}};
  dataArray_48_6_cachedata_MPORT_en_pipe_0 = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  dataArray_48_6_cachedata_MPORT_addr_pipe_0 = _RAND_2324[1:0];
  _RAND_2326 = {1{`RANDOM}};
  dataArray_48_7_cachedata_MPORT_en_pipe_0 = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  dataArray_48_7_cachedata_MPORT_addr_pipe_0 = _RAND_2327[1:0];
  _RAND_2329 = {1{`RANDOM}};
  dataArray_48_8_cachedata_MPORT_en_pipe_0 = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  dataArray_48_8_cachedata_MPORT_addr_pipe_0 = _RAND_2330[1:0];
  _RAND_2332 = {1{`RANDOM}};
  dataArray_48_9_cachedata_MPORT_en_pipe_0 = _RAND_2332[0:0];
  _RAND_2333 = {1{`RANDOM}};
  dataArray_48_9_cachedata_MPORT_addr_pipe_0 = _RAND_2333[1:0];
  _RAND_2335 = {1{`RANDOM}};
  dataArray_48_10_cachedata_MPORT_en_pipe_0 = _RAND_2335[0:0];
  _RAND_2336 = {1{`RANDOM}};
  dataArray_48_10_cachedata_MPORT_addr_pipe_0 = _RAND_2336[1:0];
  _RAND_2338 = {1{`RANDOM}};
  dataArray_48_11_cachedata_MPORT_en_pipe_0 = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  dataArray_48_11_cachedata_MPORT_addr_pipe_0 = _RAND_2339[1:0];
  _RAND_2341 = {1{`RANDOM}};
  dataArray_48_12_cachedata_MPORT_en_pipe_0 = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  dataArray_48_12_cachedata_MPORT_addr_pipe_0 = _RAND_2342[1:0];
  _RAND_2344 = {1{`RANDOM}};
  dataArray_48_13_cachedata_MPORT_en_pipe_0 = _RAND_2344[0:0];
  _RAND_2345 = {1{`RANDOM}};
  dataArray_48_13_cachedata_MPORT_addr_pipe_0 = _RAND_2345[1:0];
  _RAND_2347 = {1{`RANDOM}};
  dataArray_48_14_cachedata_MPORT_en_pipe_0 = _RAND_2347[0:0];
  _RAND_2348 = {1{`RANDOM}};
  dataArray_48_14_cachedata_MPORT_addr_pipe_0 = _RAND_2348[1:0];
  _RAND_2350 = {1{`RANDOM}};
  dataArray_48_15_cachedata_MPORT_en_pipe_0 = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  dataArray_48_15_cachedata_MPORT_addr_pipe_0 = _RAND_2351[1:0];
  _RAND_2353 = {1{`RANDOM}};
  dataArray_49_0_cachedata_MPORT_en_pipe_0 = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  dataArray_49_0_cachedata_MPORT_addr_pipe_0 = _RAND_2354[1:0];
  _RAND_2356 = {1{`RANDOM}};
  dataArray_49_1_cachedata_MPORT_en_pipe_0 = _RAND_2356[0:0];
  _RAND_2357 = {1{`RANDOM}};
  dataArray_49_1_cachedata_MPORT_addr_pipe_0 = _RAND_2357[1:0];
  _RAND_2359 = {1{`RANDOM}};
  dataArray_49_2_cachedata_MPORT_en_pipe_0 = _RAND_2359[0:0];
  _RAND_2360 = {1{`RANDOM}};
  dataArray_49_2_cachedata_MPORT_addr_pipe_0 = _RAND_2360[1:0];
  _RAND_2362 = {1{`RANDOM}};
  dataArray_49_3_cachedata_MPORT_en_pipe_0 = _RAND_2362[0:0];
  _RAND_2363 = {1{`RANDOM}};
  dataArray_49_3_cachedata_MPORT_addr_pipe_0 = _RAND_2363[1:0];
  _RAND_2365 = {1{`RANDOM}};
  dataArray_49_4_cachedata_MPORT_en_pipe_0 = _RAND_2365[0:0];
  _RAND_2366 = {1{`RANDOM}};
  dataArray_49_4_cachedata_MPORT_addr_pipe_0 = _RAND_2366[1:0];
  _RAND_2368 = {1{`RANDOM}};
  dataArray_49_5_cachedata_MPORT_en_pipe_0 = _RAND_2368[0:0];
  _RAND_2369 = {1{`RANDOM}};
  dataArray_49_5_cachedata_MPORT_addr_pipe_0 = _RAND_2369[1:0];
  _RAND_2371 = {1{`RANDOM}};
  dataArray_49_6_cachedata_MPORT_en_pipe_0 = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  dataArray_49_6_cachedata_MPORT_addr_pipe_0 = _RAND_2372[1:0];
  _RAND_2374 = {1{`RANDOM}};
  dataArray_49_7_cachedata_MPORT_en_pipe_0 = _RAND_2374[0:0];
  _RAND_2375 = {1{`RANDOM}};
  dataArray_49_7_cachedata_MPORT_addr_pipe_0 = _RAND_2375[1:0];
  _RAND_2377 = {1{`RANDOM}};
  dataArray_49_8_cachedata_MPORT_en_pipe_0 = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  dataArray_49_8_cachedata_MPORT_addr_pipe_0 = _RAND_2378[1:0];
  _RAND_2380 = {1{`RANDOM}};
  dataArray_49_9_cachedata_MPORT_en_pipe_0 = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  dataArray_49_9_cachedata_MPORT_addr_pipe_0 = _RAND_2381[1:0];
  _RAND_2383 = {1{`RANDOM}};
  dataArray_49_10_cachedata_MPORT_en_pipe_0 = _RAND_2383[0:0];
  _RAND_2384 = {1{`RANDOM}};
  dataArray_49_10_cachedata_MPORT_addr_pipe_0 = _RAND_2384[1:0];
  _RAND_2386 = {1{`RANDOM}};
  dataArray_49_11_cachedata_MPORT_en_pipe_0 = _RAND_2386[0:0];
  _RAND_2387 = {1{`RANDOM}};
  dataArray_49_11_cachedata_MPORT_addr_pipe_0 = _RAND_2387[1:0];
  _RAND_2389 = {1{`RANDOM}};
  dataArray_49_12_cachedata_MPORT_en_pipe_0 = _RAND_2389[0:0];
  _RAND_2390 = {1{`RANDOM}};
  dataArray_49_12_cachedata_MPORT_addr_pipe_0 = _RAND_2390[1:0];
  _RAND_2392 = {1{`RANDOM}};
  dataArray_49_13_cachedata_MPORT_en_pipe_0 = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  dataArray_49_13_cachedata_MPORT_addr_pipe_0 = _RAND_2393[1:0];
  _RAND_2395 = {1{`RANDOM}};
  dataArray_49_14_cachedata_MPORT_en_pipe_0 = _RAND_2395[0:0];
  _RAND_2396 = {1{`RANDOM}};
  dataArray_49_14_cachedata_MPORT_addr_pipe_0 = _RAND_2396[1:0];
  _RAND_2398 = {1{`RANDOM}};
  dataArray_49_15_cachedata_MPORT_en_pipe_0 = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  dataArray_49_15_cachedata_MPORT_addr_pipe_0 = _RAND_2399[1:0];
  _RAND_2401 = {1{`RANDOM}};
  dataArray_50_0_cachedata_MPORT_en_pipe_0 = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  dataArray_50_0_cachedata_MPORT_addr_pipe_0 = _RAND_2402[1:0];
  _RAND_2404 = {1{`RANDOM}};
  dataArray_50_1_cachedata_MPORT_en_pipe_0 = _RAND_2404[0:0];
  _RAND_2405 = {1{`RANDOM}};
  dataArray_50_1_cachedata_MPORT_addr_pipe_0 = _RAND_2405[1:0];
  _RAND_2407 = {1{`RANDOM}};
  dataArray_50_2_cachedata_MPORT_en_pipe_0 = _RAND_2407[0:0];
  _RAND_2408 = {1{`RANDOM}};
  dataArray_50_2_cachedata_MPORT_addr_pipe_0 = _RAND_2408[1:0];
  _RAND_2410 = {1{`RANDOM}};
  dataArray_50_3_cachedata_MPORT_en_pipe_0 = _RAND_2410[0:0];
  _RAND_2411 = {1{`RANDOM}};
  dataArray_50_3_cachedata_MPORT_addr_pipe_0 = _RAND_2411[1:0];
  _RAND_2413 = {1{`RANDOM}};
  dataArray_50_4_cachedata_MPORT_en_pipe_0 = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  dataArray_50_4_cachedata_MPORT_addr_pipe_0 = _RAND_2414[1:0];
  _RAND_2416 = {1{`RANDOM}};
  dataArray_50_5_cachedata_MPORT_en_pipe_0 = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  dataArray_50_5_cachedata_MPORT_addr_pipe_0 = _RAND_2417[1:0];
  _RAND_2419 = {1{`RANDOM}};
  dataArray_50_6_cachedata_MPORT_en_pipe_0 = _RAND_2419[0:0];
  _RAND_2420 = {1{`RANDOM}};
  dataArray_50_6_cachedata_MPORT_addr_pipe_0 = _RAND_2420[1:0];
  _RAND_2422 = {1{`RANDOM}};
  dataArray_50_7_cachedata_MPORT_en_pipe_0 = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  dataArray_50_7_cachedata_MPORT_addr_pipe_0 = _RAND_2423[1:0];
  _RAND_2425 = {1{`RANDOM}};
  dataArray_50_8_cachedata_MPORT_en_pipe_0 = _RAND_2425[0:0];
  _RAND_2426 = {1{`RANDOM}};
  dataArray_50_8_cachedata_MPORT_addr_pipe_0 = _RAND_2426[1:0];
  _RAND_2428 = {1{`RANDOM}};
  dataArray_50_9_cachedata_MPORT_en_pipe_0 = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  dataArray_50_9_cachedata_MPORT_addr_pipe_0 = _RAND_2429[1:0];
  _RAND_2431 = {1{`RANDOM}};
  dataArray_50_10_cachedata_MPORT_en_pipe_0 = _RAND_2431[0:0];
  _RAND_2432 = {1{`RANDOM}};
  dataArray_50_10_cachedata_MPORT_addr_pipe_0 = _RAND_2432[1:0];
  _RAND_2434 = {1{`RANDOM}};
  dataArray_50_11_cachedata_MPORT_en_pipe_0 = _RAND_2434[0:0];
  _RAND_2435 = {1{`RANDOM}};
  dataArray_50_11_cachedata_MPORT_addr_pipe_0 = _RAND_2435[1:0];
  _RAND_2437 = {1{`RANDOM}};
  dataArray_50_12_cachedata_MPORT_en_pipe_0 = _RAND_2437[0:0];
  _RAND_2438 = {1{`RANDOM}};
  dataArray_50_12_cachedata_MPORT_addr_pipe_0 = _RAND_2438[1:0];
  _RAND_2440 = {1{`RANDOM}};
  dataArray_50_13_cachedata_MPORT_en_pipe_0 = _RAND_2440[0:0];
  _RAND_2441 = {1{`RANDOM}};
  dataArray_50_13_cachedata_MPORT_addr_pipe_0 = _RAND_2441[1:0];
  _RAND_2443 = {1{`RANDOM}};
  dataArray_50_14_cachedata_MPORT_en_pipe_0 = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  dataArray_50_14_cachedata_MPORT_addr_pipe_0 = _RAND_2444[1:0];
  _RAND_2446 = {1{`RANDOM}};
  dataArray_50_15_cachedata_MPORT_en_pipe_0 = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  dataArray_50_15_cachedata_MPORT_addr_pipe_0 = _RAND_2447[1:0];
  _RAND_2449 = {1{`RANDOM}};
  dataArray_51_0_cachedata_MPORT_en_pipe_0 = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  dataArray_51_0_cachedata_MPORT_addr_pipe_0 = _RAND_2450[1:0];
  _RAND_2452 = {1{`RANDOM}};
  dataArray_51_1_cachedata_MPORT_en_pipe_0 = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  dataArray_51_1_cachedata_MPORT_addr_pipe_0 = _RAND_2453[1:0];
  _RAND_2455 = {1{`RANDOM}};
  dataArray_51_2_cachedata_MPORT_en_pipe_0 = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  dataArray_51_2_cachedata_MPORT_addr_pipe_0 = _RAND_2456[1:0];
  _RAND_2458 = {1{`RANDOM}};
  dataArray_51_3_cachedata_MPORT_en_pipe_0 = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  dataArray_51_3_cachedata_MPORT_addr_pipe_0 = _RAND_2459[1:0];
  _RAND_2461 = {1{`RANDOM}};
  dataArray_51_4_cachedata_MPORT_en_pipe_0 = _RAND_2461[0:0];
  _RAND_2462 = {1{`RANDOM}};
  dataArray_51_4_cachedata_MPORT_addr_pipe_0 = _RAND_2462[1:0];
  _RAND_2464 = {1{`RANDOM}};
  dataArray_51_5_cachedata_MPORT_en_pipe_0 = _RAND_2464[0:0];
  _RAND_2465 = {1{`RANDOM}};
  dataArray_51_5_cachedata_MPORT_addr_pipe_0 = _RAND_2465[1:0];
  _RAND_2467 = {1{`RANDOM}};
  dataArray_51_6_cachedata_MPORT_en_pipe_0 = _RAND_2467[0:0];
  _RAND_2468 = {1{`RANDOM}};
  dataArray_51_6_cachedata_MPORT_addr_pipe_0 = _RAND_2468[1:0];
  _RAND_2470 = {1{`RANDOM}};
  dataArray_51_7_cachedata_MPORT_en_pipe_0 = _RAND_2470[0:0];
  _RAND_2471 = {1{`RANDOM}};
  dataArray_51_7_cachedata_MPORT_addr_pipe_0 = _RAND_2471[1:0];
  _RAND_2473 = {1{`RANDOM}};
  dataArray_51_8_cachedata_MPORT_en_pipe_0 = _RAND_2473[0:0];
  _RAND_2474 = {1{`RANDOM}};
  dataArray_51_8_cachedata_MPORT_addr_pipe_0 = _RAND_2474[1:0];
  _RAND_2476 = {1{`RANDOM}};
  dataArray_51_9_cachedata_MPORT_en_pipe_0 = _RAND_2476[0:0];
  _RAND_2477 = {1{`RANDOM}};
  dataArray_51_9_cachedata_MPORT_addr_pipe_0 = _RAND_2477[1:0];
  _RAND_2479 = {1{`RANDOM}};
  dataArray_51_10_cachedata_MPORT_en_pipe_0 = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  dataArray_51_10_cachedata_MPORT_addr_pipe_0 = _RAND_2480[1:0];
  _RAND_2482 = {1{`RANDOM}};
  dataArray_51_11_cachedata_MPORT_en_pipe_0 = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  dataArray_51_11_cachedata_MPORT_addr_pipe_0 = _RAND_2483[1:0];
  _RAND_2485 = {1{`RANDOM}};
  dataArray_51_12_cachedata_MPORT_en_pipe_0 = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  dataArray_51_12_cachedata_MPORT_addr_pipe_0 = _RAND_2486[1:0];
  _RAND_2488 = {1{`RANDOM}};
  dataArray_51_13_cachedata_MPORT_en_pipe_0 = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  dataArray_51_13_cachedata_MPORT_addr_pipe_0 = _RAND_2489[1:0];
  _RAND_2491 = {1{`RANDOM}};
  dataArray_51_14_cachedata_MPORT_en_pipe_0 = _RAND_2491[0:0];
  _RAND_2492 = {1{`RANDOM}};
  dataArray_51_14_cachedata_MPORT_addr_pipe_0 = _RAND_2492[1:0];
  _RAND_2494 = {1{`RANDOM}};
  dataArray_51_15_cachedata_MPORT_en_pipe_0 = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  dataArray_51_15_cachedata_MPORT_addr_pipe_0 = _RAND_2495[1:0];
  _RAND_2497 = {1{`RANDOM}};
  dataArray_52_0_cachedata_MPORT_en_pipe_0 = _RAND_2497[0:0];
  _RAND_2498 = {1{`RANDOM}};
  dataArray_52_0_cachedata_MPORT_addr_pipe_0 = _RAND_2498[1:0];
  _RAND_2500 = {1{`RANDOM}};
  dataArray_52_1_cachedata_MPORT_en_pipe_0 = _RAND_2500[0:0];
  _RAND_2501 = {1{`RANDOM}};
  dataArray_52_1_cachedata_MPORT_addr_pipe_0 = _RAND_2501[1:0];
  _RAND_2503 = {1{`RANDOM}};
  dataArray_52_2_cachedata_MPORT_en_pipe_0 = _RAND_2503[0:0];
  _RAND_2504 = {1{`RANDOM}};
  dataArray_52_2_cachedata_MPORT_addr_pipe_0 = _RAND_2504[1:0];
  _RAND_2506 = {1{`RANDOM}};
  dataArray_52_3_cachedata_MPORT_en_pipe_0 = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  dataArray_52_3_cachedata_MPORT_addr_pipe_0 = _RAND_2507[1:0];
  _RAND_2509 = {1{`RANDOM}};
  dataArray_52_4_cachedata_MPORT_en_pipe_0 = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  dataArray_52_4_cachedata_MPORT_addr_pipe_0 = _RAND_2510[1:0];
  _RAND_2512 = {1{`RANDOM}};
  dataArray_52_5_cachedata_MPORT_en_pipe_0 = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  dataArray_52_5_cachedata_MPORT_addr_pipe_0 = _RAND_2513[1:0];
  _RAND_2515 = {1{`RANDOM}};
  dataArray_52_6_cachedata_MPORT_en_pipe_0 = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  dataArray_52_6_cachedata_MPORT_addr_pipe_0 = _RAND_2516[1:0];
  _RAND_2518 = {1{`RANDOM}};
  dataArray_52_7_cachedata_MPORT_en_pipe_0 = _RAND_2518[0:0];
  _RAND_2519 = {1{`RANDOM}};
  dataArray_52_7_cachedata_MPORT_addr_pipe_0 = _RAND_2519[1:0];
  _RAND_2521 = {1{`RANDOM}};
  dataArray_52_8_cachedata_MPORT_en_pipe_0 = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  dataArray_52_8_cachedata_MPORT_addr_pipe_0 = _RAND_2522[1:0];
  _RAND_2524 = {1{`RANDOM}};
  dataArray_52_9_cachedata_MPORT_en_pipe_0 = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  dataArray_52_9_cachedata_MPORT_addr_pipe_0 = _RAND_2525[1:0];
  _RAND_2527 = {1{`RANDOM}};
  dataArray_52_10_cachedata_MPORT_en_pipe_0 = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  dataArray_52_10_cachedata_MPORT_addr_pipe_0 = _RAND_2528[1:0];
  _RAND_2530 = {1{`RANDOM}};
  dataArray_52_11_cachedata_MPORT_en_pipe_0 = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  dataArray_52_11_cachedata_MPORT_addr_pipe_0 = _RAND_2531[1:0];
  _RAND_2533 = {1{`RANDOM}};
  dataArray_52_12_cachedata_MPORT_en_pipe_0 = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  dataArray_52_12_cachedata_MPORT_addr_pipe_0 = _RAND_2534[1:0];
  _RAND_2536 = {1{`RANDOM}};
  dataArray_52_13_cachedata_MPORT_en_pipe_0 = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  dataArray_52_13_cachedata_MPORT_addr_pipe_0 = _RAND_2537[1:0];
  _RAND_2539 = {1{`RANDOM}};
  dataArray_52_14_cachedata_MPORT_en_pipe_0 = _RAND_2539[0:0];
  _RAND_2540 = {1{`RANDOM}};
  dataArray_52_14_cachedata_MPORT_addr_pipe_0 = _RAND_2540[1:0];
  _RAND_2542 = {1{`RANDOM}};
  dataArray_52_15_cachedata_MPORT_en_pipe_0 = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  dataArray_52_15_cachedata_MPORT_addr_pipe_0 = _RAND_2543[1:0];
  _RAND_2545 = {1{`RANDOM}};
  dataArray_53_0_cachedata_MPORT_en_pipe_0 = _RAND_2545[0:0];
  _RAND_2546 = {1{`RANDOM}};
  dataArray_53_0_cachedata_MPORT_addr_pipe_0 = _RAND_2546[1:0];
  _RAND_2548 = {1{`RANDOM}};
  dataArray_53_1_cachedata_MPORT_en_pipe_0 = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  dataArray_53_1_cachedata_MPORT_addr_pipe_0 = _RAND_2549[1:0];
  _RAND_2551 = {1{`RANDOM}};
  dataArray_53_2_cachedata_MPORT_en_pipe_0 = _RAND_2551[0:0];
  _RAND_2552 = {1{`RANDOM}};
  dataArray_53_2_cachedata_MPORT_addr_pipe_0 = _RAND_2552[1:0];
  _RAND_2554 = {1{`RANDOM}};
  dataArray_53_3_cachedata_MPORT_en_pipe_0 = _RAND_2554[0:0];
  _RAND_2555 = {1{`RANDOM}};
  dataArray_53_3_cachedata_MPORT_addr_pipe_0 = _RAND_2555[1:0];
  _RAND_2557 = {1{`RANDOM}};
  dataArray_53_4_cachedata_MPORT_en_pipe_0 = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  dataArray_53_4_cachedata_MPORT_addr_pipe_0 = _RAND_2558[1:0];
  _RAND_2560 = {1{`RANDOM}};
  dataArray_53_5_cachedata_MPORT_en_pipe_0 = _RAND_2560[0:0];
  _RAND_2561 = {1{`RANDOM}};
  dataArray_53_5_cachedata_MPORT_addr_pipe_0 = _RAND_2561[1:0];
  _RAND_2563 = {1{`RANDOM}};
  dataArray_53_6_cachedata_MPORT_en_pipe_0 = _RAND_2563[0:0];
  _RAND_2564 = {1{`RANDOM}};
  dataArray_53_6_cachedata_MPORT_addr_pipe_0 = _RAND_2564[1:0];
  _RAND_2566 = {1{`RANDOM}};
  dataArray_53_7_cachedata_MPORT_en_pipe_0 = _RAND_2566[0:0];
  _RAND_2567 = {1{`RANDOM}};
  dataArray_53_7_cachedata_MPORT_addr_pipe_0 = _RAND_2567[1:0];
  _RAND_2569 = {1{`RANDOM}};
  dataArray_53_8_cachedata_MPORT_en_pipe_0 = _RAND_2569[0:0];
  _RAND_2570 = {1{`RANDOM}};
  dataArray_53_8_cachedata_MPORT_addr_pipe_0 = _RAND_2570[1:0];
  _RAND_2572 = {1{`RANDOM}};
  dataArray_53_9_cachedata_MPORT_en_pipe_0 = _RAND_2572[0:0];
  _RAND_2573 = {1{`RANDOM}};
  dataArray_53_9_cachedata_MPORT_addr_pipe_0 = _RAND_2573[1:0];
  _RAND_2575 = {1{`RANDOM}};
  dataArray_53_10_cachedata_MPORT_en_pipe_0 = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  dataArray_53_10_cachedata_MPORT_addr_pipe_0 = _RAND_2576[1:0];
  _RAND_2578 = {1{`RANDOM}};
  dataArray_53_11_cachedata_MPORT_en_pipe_0 = _RAND_2578[0:0];
  _RAND_2579 = {1{`RANDOM}};
  dataArray_53_11_cachedata_MPORT_addr_pipe_0 = _RAND_2579[1:0];
  _RAND_2581 = {1{`RANDOM}};
  dataArray_53_12_cachedata_MPORT_en_pipe_0 = _RAND_2581[0:0];
  _RAND_2582 = {1{`RANDOM}};
  dataArray_53_12_cachedata_MPORT_addr_pipe_0 = _RAND_2582[1:0];
  _RAND_2584 = {1{`RANDOM}};
  dataArray_53_13_cachedata_MPORT_en_pipe_0 = _RAND_2584[0:0];
  _RAND_2585 = {1{`RANDOM}};
  dataArray_53_13_cachedata_MPORT_addr_pipe_0 = _RAND_2585[1:0];
  _RAND_2587 = {1{`RANDOM}};
  dataArray_53_14_cachedata_MPORT_en_pipe_0 = _RAND_2587[0:0];
  _RAND_2588 = {1{`RANDOM}};
  dataArray_53_14_cachedata_MPORT_addr_pipe_0 = _RAND_2588[1:0];
  _RAND_2590 = {1{`RANDOM}};
  dataArray_53_15_cachedata_MPORT_en_pipe_0 = _RAND_2590[0:0];
  _RAND_2591 = {1{`RANDOM}};
  dataArray_53_15_cachedata_MPORT_addr_pipe_0 = _RAND_2591[1:0];
  _RAND_2593 = {1{`RANDOM}};
  dataArray_54_0_cachedata_MPORT_en_pipe_0 = _RAND_2593[0:0];
  _RAND_2594 = {1{`RANDOM}};
  dataArray_54_0_cachedata_MPORT_addr_pipe_0 = _RAND_2594[1:0];
  _RAND_2596 = {1{`RANDOM}};
  dataArray_54_1_cachedata_MPORT_en_pipe_0 = _RAND_2596[0:0];
  _RAND_2597 = {1{`RANDOM}};
  dataArray_54_1_cachedata_MPORT_addr_pipe_0 = _RAND_2597[1:0];
  _RAND_2599 = {1{`RANDOM}};
  dataArray_54_2_cachedata_MPORT_en_pipe_0 = _RAND_2599[0:0];
  _RAND_2600 = {1{`RANDOM}};
  dataArray_54_2_cachedata_MPORT_addr_pipe_0 = _RAND_2600[1:0];
  _RAND_2602 = {1{`RANDOM}};
  dataArray_54_3_cachedata_MPORT_en_pipe_0 = _RAND_2602[0:0];
  _RAND_2603 = {1{`RANDOM}};
  dataArray_54_3_cachedata_MPORT_addr_pipe_0 = _RAND_2603[1:0];
  _RAND_2605 = {1{`RANDOM}};
  dataArray_54_4_cachedata_MPORT_en_pipe_0 = _RAND_2605[0:0];
  _RAND_2606 = {1{`RANDOM}};
  dataArray_54_4_cachedata_MPORT_addr_pipe_0 = _RAND_2606[1:0];
  _RAND_2608 = {1{`RANDOM}};
  dataArray_54_5_cachedata_MPORT_en_pipe_0 = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  dataArray_54_5_cachedata_MPORT_addr_pipe_0 = _RAND_2609[1:0];
  _RAND_2611 = {1{`RANDOM}};
  dataArray_54_6_cachedata_MPORT_en_pipe_0 = _RAND_2611[0:0];
  _RAND_2612 = {1{`RANDOM}};
  dataArray_54_6_cachedata_MPORT_addr_pipe_0 = _RAND_2612[1:0];
  _RAND_2614 = {1{`RANDOM}};
  dataArray_54_7_cachedata_MPORT_en_pipe_0 = _RAND_2614[0:0];
  _RAND_2615 = {1{`RANDOM}};
  dataArray_54_7_cachedata_MPORT_addr_pipe_0 = _RAND_2615[1:0];
  _RAND_2617 = {1{`RANDOM}};
  dataArray_54_8_cachedata_MPORT_en_pipe_0 = _RAND_2617[0:0];
  _RAND_2618 = {1{`RANDOM}};
  dataArray_54_8_cachedata_MPORT_addr_pipe_0 = _RAND_2618[1:0];
  _RAND_2620 = {1{`RANDOM}};
  dataArray_54_9_cachedata_MPORT_en_pipe_0 = _RAND_2620[0:0];
  _RAND_2621 = {1{`RANDOM}};
  dataArray_54_9_cachedata_MPORT_addr_pipe_0 = _RAND_2621[1:0];
  _RAND_2623 = {1{`RANDOM}};
  dataArray_54_10_cachedata_MPORT_en_pipe_0 = _RAND_2623[0:0];
  _RAND_2624 = {1{`RANDOM}};
  dataArray_54_10_cachedata_MPORT_addr_pipe_0 = _RAND_2624[1:0];
  _RAND_2626 = {1{`RANDOM}};
  dataArray_54_11_cachedata_MPORT_en_pipe_0 = _RAND_2626[0:0];
  _RAND_2627 = {1{`RANDOM}};
  dataArray_54_11_cachedata_MPORT_addr_pipe_0 = _RAND_2627[1:0];
  _RAND_2629 = {1{`RANDOM}};
  dataArray_54_12_cachedata_MPORT_en_pipe_0 = _RAND_2629[0:0];
  _RAND_2630 = {1{`RANDOM}};
  dataArray_54_12_cachedata_MPORT_addr_pipe_0 = _RAND_2630[1:0];
  _RAND_2632 = {1{`RANDOM}};
  dataArray_54_13_cachedata_MPORT_en_pipe_0 = _RAND_2632[0:0];
  _RAND_2633 = {1{`RANDOM}};
  dataArray_54_13_cachedata_MPORT_addr_pipe_0 = _RAND_2633[1:0];
  _RAND_2635 = {1{`RANDOM}};
  dataArray_54_14_cachedata_MPORT_en_pipe_0 = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  dataArray_54_14_cachedata_MPORT_addr_pipe_0 = _RAND_2636[1:0];
  _RAND_2638 = {1{`RANDOM}};
  dataArray_54_15_cachedata_MPORT_en_pipe_0 = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  dataArray_54_15_cachedata_MPORT_addr_pipe_0 = _RAND_2639[1:0];
  _RAND_2641 = {1{`RANDOM}};
  dataArray_55_0_cachedata_MPORT_en_pipe_0 = _RAND_2641[0:0];
  _RAND_2642 = {1{`RANDOM}};
  dataArray_55_0_cachedata_MPORT_addr_pipe_0 = _RAND_2642[1:0];
  _RAND_2644 = {1{`RANDOM}};
  dataArray_55_1_cachedata_MPORT_en_pipe_0 = _RAND_2644[0:0];
  _RAND_2645 = {1{`RANDOM}};
  dataArray_55_1_cachedata_MPORT_addr_pipe_0 = _RAND_2645[1:0];
  _RAND_2647 = {1{`RANDOM}};
  dataArray_55_2_cachedata_MPORT_en_pipe_0 = _RAND_2647[0:0];
  _RAND_2648 = {1{`RANDOM}};
  dataArray_55_2_cachedata_MPORT_addr_pipe_0 = _RAND_2648[1:0];
  _RAND_2650 = {1{`RANDOM}};
  dataArray_55_3_cachedata_MPORT_en_pipe_0 = _RAND_2650[0:0];
  _RAND_2651 = {1{`RANDOM}};
  dataArray_55_3_cachedata_MPORT_addr_pipe_0 = _RAND_2651[1:0];
  _RAND_2653 = {1{`RANDOM}};
  dataArray_55_4_cachedata_MPORT_en_pipe_0 = _RAND_2653[0:0];
  _RAND_2654 = {1{`RANDOM}};
  dataArray_55_4_cachedata_MPORT_addr_pipe_0 = _RAND_2654[1:0];
  _RAND_2656 = {1{`RANDOM}};
  dataArray_55_5_cachedata_MPORT_en_pipe_0 = _RAND_2656[0:0];
  _RAND_2657 = {1{`RANDOM}};
  dataArray_55_5_cachedata_MPORT_addr_pipe_0 = _RAND_2657[1:0];
  _RAND_2659 = {1{`RANDOM}};
  dataArray_55_6_cachedata_MPORT_en_pipe_0 = _RAND_2659[0:0];
  _RAND_2660 = {1{`RANDOM}};
  dataArray_55_6_cachedata_MPORT_addr_pipe_0 = _RAND_2660[1:0];
  _RAND_2662 = {1{`RANDOM}};
  dataArray_55_7_cachedata_MPORT_en_pipe_0 = _RAND_2662[0:0];
  _RAND_2663 = {1{`RANDOM}};
  dataArray_55_7_cachedata_MPORT_addr_pipe_0 = _RAND_2663[1:0];
  _RAND_2665 = {1{`RANDOM}};
  dataArray_55_8_cachedata_MPORT_en_pipe_0 = _RAND_2665[0:0];
  _RAND_2666 = {1{`RANDOM}};
  dataArray_55_8_cachedata_MPORT_addr_pipe_0 = _RAND_2666[1:0];
  _RAND_2668 = {1{`RANDOM}};
  dataArray_55_9_cachedata_MPORT_en_pipe_0 = _RAND_2668[0:0];
  _RAND_2669 = {1{`RANDOM}};
  dataArray_55_9_cachedata_MPORT_addr_pipe_0 = _RAND_2669[1:0];
  _RAND_2671 = {1{`RANDOM}};
  dataArray_55_10_cachedata_MPORT_en_pipe_0 = _RAND_2671[0:0];
  _RAND_2672 = {1{`RANDOM}};
  dataArray_55_10_cachedata_MPORT_addr_pipe_0 = _RAND_2672[1:0];
  _RAND_2674 = {1{`RANDOM}};
  dataArray_55_11_cachedata_MPORT_en_pipe_0 = _RAND_2674[0:0];
  _RAND_2675 = {1{`RANDOM}};
  dataArray_55_11_cachedata_MPORT_addr_pipe_0 = _RAND_2675[1:0];
  _RAND_2677 = {1{`RANDOM}};
  dataArray_55_12_cachedata_MPORT_en_pipe_0 = _RAND_2677[0:0];
  _RAND_2678 = {1{`RANDOM}};
  dataArray_55_12_cachedata_MPORT_addr_pipe_0 = _RAND_2678[1:0];
  _RAND_2680 = {1{`RANDOM}};
  dataArray_55_13_cachedata_MPORT_en_pipe_0 = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  dataArray_55_13_cachedata_MPORT_addr_pipe_0 = _RAND_2681[1:0];
  _RAND_2683 = {1{`RANDOM}};
  dataArray_55_14_cachedata_MPORT_en_pipe_0 = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  dataArray_55_14_cachedata_MPORT_addr_pipe_0 = _RAND_2684[1:0];
  _RAND_2686 = {1{`RANDOM}};
  dataArray_55_15_cachedata_MPORT_en_pipe_0 = _RAND_2686[0:0];
  _RAND_2687 = {1{`RANDOM}};
  dataArray_55_15_cachedata_MPORT_addr_pipe_0 = _RAND_2687[1:0];
  _RAND_2689 = {1{`RANDOM}};
  dataArray_56_0_cachedata_MPORT_en_pipe_0 = _RAND_2689[0:0];
  _RAND_2690 = {1{`RANDOM}};
  dataArray_56_0_cachedata_MPORT_addr_pipe_0 = _RAND_2690[1:0];
  _RAND_2692 = {1{`RANDOM}};
  dataArray_56_1_cachedata_MPORT_en_pipe_0 = _RAND_2692[0:0];
  _RAND_2693 = {1{`RANDOM}};
  dataArray_56_1_cachedata_MPORT_addr_pipe_0 = _RAND_2693[1:0];
  _RAND_2695 = {1{`RANDOM}};
  dataArray_56_2_cachedata_MPORT_en_pipe_0 = _RAND_2695[0:0];
  _RAND_2696 = {1{`RANDOM}};
  dataArray_56_2_cachedata_MPORT_addr_pipe_0 = _RAND_2696[1:0];
  _RAND_2698 = {1{`RANDOM}};
  dataArray_56_3_cachedata_MPORT_en_pipe_0 = _RAND_2698[0:0];
  _RAND_2699 = {1{`RANDOM}};
  dataArray_56_3_cachedata_MPORT_addr_pipe_0 = _RAND_2699[1:0];
  _RAND_2701 = {1{`RANDOM}};
  dataArray_56_4_cachedata_MPORT_en_pipe_0 = _RAND_2701[0:0];
  _RAND_2702 = {1{`RANDOM}};
  dataArray_56_4_cachedata_MPORT_addr_pipe_0 = _RAND_2702[1:0];
  _RAND_2704 = {1{`RANDOM}};
  dataArray_56_5_cachedata_MPORT_en_pipe_0 = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  dataArray_56_5_cachedata_MPORT_addr_pipe_0 = _RAND_2705[1:0];
  _RAND_2707 = {1{`RANDOM}};
  dataArray_56_6_cachedata_MPORT_en_pipe_0 = _RAND_2707[0:0];
  _RAND_2708 = {1{`RANDOM}};
  dataArray_56_6_cachedata_MPORT_addr_pipe_0 = _RAND_2708[1:0];
  _RAND_2710 = {1{`RANDOM}};
  dataArray_56_7_cachedata_MPORT_en_pipe_0 = _RAND_2710[0:0];
  _RAND_2711 = {1{`RANDOM}};
  dataArray_56_7_cachedata_MPORT_addr_pipe_0 = _RAND_2711[1:0];
  _RAND_2713 = {1{`RANDOM}};
  dataArray_56_8_cachedata_MPORT_en_pipe_0 = _RAND_2713[0:0];
  _RAND_2714 = {1{`RANDOM}};
  dataArray_56_8_cachedata_MPORT_addr_pipe_0 = _RAND_2714[1:0];
  _RAND_2716 = {1{`RANDOM}};
  dataArray_56_9_cachedata_MPORT_en_pipe_0 = _RAND_2716[0:0];
  _RAND_2717 = {1{`RANDOM}};
  dataArray_56_9_cachedata_MPORT_addr_pipe_0 = _RAND_2717[1:0];
  _RAND_2719 = {1{`RANDOM}};
  dataArray_56_10_cachedata_MPORT_en_pipe_0 = _RAND_2719[0:0];
  _RAND_2720 = {1{`RANDOM}};
  dataArray_56_10_cachedata_MPORT_addr_pipe_0 = _RAND_2720[1:0];
  _RAND_2722 = {1{`RANDOM}};
  dataArray_56_11_cachedata_MPORT_en_pipe_0 = _RAND_2722[0:0];
  _RAND_2723 = {1{`RANDOM}};
  dataArray_56_11_cachedata_MPORT_addr_pipe_0 = _RAND_2723[1:0];
  _RAND_2725 = {1{`RANDOM}};
  dataArray_56_12_cachedata_MPORT_en_pipe_0 = _RAND_2725[0:0];
  _RAND_2726 = {1{`RANDOM}};
  dataArray_56_12_cachedata_MPORT_addr_pipe_0 = _RAND_2726[1:0];
  _RAND_2728 = {1{`RANDOM}};
  dataArray_56_13_cachedata_MPORT_en_pipe_0 = _RAND_2728[0:0];
  _RAND_2729 = {1{`RANDOM}};
  dataArray_56_13_cachedata_MPORT_addr_pipe_0 = _RAND_2729[1:0];
  _RAND_2731 = {1{`RANDOM}};
  dataArray_56_14_cachedata_MPORT_en_pipe_0 = _RAND_2731[0:0];
  _RAND_2732 = {1{`RANDOM}};
  dataArray_56_14_cachedata_MPORT_addr_pipe_0 = _RAND_2732[1:0];
  _RAND_2734 = {1{`RANDOM}};
  dataArray_56_15_cachedata_MPORT_en_pipe_0 = _RAND_2734[0:0];
  _RAND_2735 = {1{`RANDOM}};
  dataArray_56_15_cachedata_MPORT_addr_pipe_0 = _RAND_2735[1:0];
  _RAND_2737 = {1{`RANDOM}};
  dataArray_57_0_cachedata_MPORT_en_pipe_0 = _RAND_2737[0:0];
  _RAND_2738 = {1{`RANDOM}};
  dataArray_57_0_cachedata_MPORT_addr_pipe_0 = _RAND_2738[1:0];
  _RAND_2740 = {1{`RANDOM}};
  dataArray_57_1_cachedata_MPORT_en_pipe_0 = _RAND_2740[0:0];
  _RAND_2741 = {1{`RANDOM}};
  dataArray_57_1_cachedata_MPORT_addr_pipe_0 = _RAND_2741[1:0];
  _RAND_2743 = {1{`RANDOM}};
  dataArray_57_2_cachedata_MPORT_en_pipe_0 = _RAND_2743[0:0];
  _RAND_2744 = {1{`RANDOM}};
  dataArray_57_2_cachedata_MPORT_addr_pipe_0 = _RAND_2744[1:0];
  _RAND_2746 = {1{`RANDOM}};
  dataArray_57_3_cachedata_MPORT_en_pipe_0 = _RAND_2746[0:0];
  _RAND_2747 = {1{`RANDOM}};
  dataArray_57_3_cachedata_MPORT_addr_pipe_0 = _RAND_2747[1:0];
  _RAND_2749 = {1{`RANDOM}};
  dataArray_57_4_cachedata_MPORT_en_pipe_0 = _RAND_2749[0:0];
  _RAND_2750 = {1{`RANDOM}};
  dataArray_57_4_cachedata_MPORT_addr_pipe_0 = _RAND_2750[1:0];
  _RAND_2752 = {1{`RANDOM}};
  dataArray_57_5_cachedata_MPORT_en_pipe_0 = _RAND_2752[0:0];
  _RAND_2753 = {1{`RANDOM}};
  dataArray_57_5_cachedata_MPORT_addr_pipe_0 = _RAND_2753[1:0];
  _RAND_2755 = {1{`RANDOM}};
  dataArray_57_6_cachedata_MPORT_en_pipe_0 = _RAND_2755[0:0];
  _RAND_2756 = {1{`RANDOM}};
  dataArray_57_6_cachedata_MPORT_addr_pipe_0 = _RAND_2756[1:0];
  _RAND_2758 = {1{`RANDOM}};
  dataArray_57_7_cachedata_MPORT_en_pipe_0 = _RAND_2758[0:0];
  _RAND_2759 = {1{`RANDOM}};
  dataArray_57_7_cachedata_MPORT_addr_pipe_0 = _RAND_2759[1:0];
  _RAND_2761 = {1{`RANDOM}};
  dataArray_57_8_cachedata_MPORT_en_pipe_0 = _RAND_2761[0:0];
  _RAND_2762 = {1{`RANDOM}};
  dataArray_57_8_cachedata_MPORT_addr_pipe_0 = _RAND_2762[1:0];
  _RAND_2764 = {1{`RANDOM}};
  dataArray_57_9_cachedata_MPORT_en_pipe_0 = _RAND_2764[0:0];
  _RAND_2765 = {1{`RANDOM}};
  dataArray_57_9_cachedata_MPORT_addr_pipe_0 = _RAND_2765[1:0];
  _RAND_2767 = {1{`RANDOM}};
  dataArray_57_10_cachedata_MPORT_en_pipe_0 = _RAND_2767[0:0];
  _RAND_2768 = {1{`RANDOM}};
  dataArray_57_10_cachedata_MPORT_addr_pipe_0 = _RAND_2768[1:0];
  _RAND_2770 = {1{`RANDOM}};
  dataArray_57_11_cachedata_MPORT_en_pipe_0 = _RAND_2770[0:0];
  _RAND_2771 = {1{`RANDOM}};
  dataArray_57_11_cachedata_MPORT_addr_pipe_0 = _RAND_2771[1:0];
  _RAND_2773 = {1{`RANDOM}};
  dataArray_57_12_cachedata_MPORT_en_pipe_0 = _RAND_2773[0:0];
  _RAND_2774 = {1{`RANDOM}};
  dataArray_57_12_cachedata_MPORT_addr_pipe_0 = _RAND_2774[1:0];
  _RAND_2776 = {1{`RANDOM}};
  dataArray_57_13_cachedata_MPORT_en_pipe_0 = _RAND_2776[0:0];
  _RAND_2777 = {1{`RANDOM}};
  dataArray_57_13_cachedata_MPORT_addr_pipe_0 = _RAND_2777[1:0];
  _RAND_2779 = {1{`RANDOM}};
  dataArray_57_14_cachedata_MPORT_en_pipe_0 = _RAND_2779[0:0];
  _RAND_2780 = {1{`RANDOM}};
  dataArray_57_14_cachedata_MPORT_addr_pipe_0 = _RAND_2780[1:0];
  _RAND_2782 = {1{`RANDOM}};
  dataArray_57_15_cachedata_MPORT_en_pipe_0 = _RAND_2782[0:0];
  _RAND_2783 = {1{`RANDOM}};
  dataArray_57_15_cachedata_MPORT_addr_pipe_0 = _RAND_2783[1:0];
  _RAND_2785 = {1{`RANDOM}};
  dataArray_58_0_cachedata_MPORT_en_pipe_0 = _RAND_2785[0:0];
  _RAND_2786 = {1{`RANDOM}};
  dataArray_58_0_cachedata_MPORT_addr_pipe_0 = _RAND_2786[1:0];
  _RAND_2788 = {1{`RANDOM}};
  dataArray_58_1_cachedata_MPORT_en_pipe_0 = _RAND_2788[0:0];
  _RAND_2789 = {1{`RANDOM}};
  dataArray_58_1_cachedata_MPORT_addr_pipe_0 = _RAND_2789[1:0];
  _RAND_2791 = {1{`RANDOM}};
  dataArray_58_2_cachedata_MPORT_en_pipe_0 = _RAND_2791[0:0];
  _RAND_2792 = {1{`RANDOM}};
  dataArray_58_2_cachedata_MPORT_addr_pipe_0 = _RAND_2792[1:0];
  _RAND_2794 = {1{`RANDOM}};
  dataArray_58_3_cachedata_MPORT_en_pipe_0 = _RAND_2794[0:0];
  _RAND_2795 = {1{`RANDOM}};
  dataArray_58_3_cachedata_MPORT_addr_pipe_0 = _RAND_2795[1:0];
  _RAND_2797 = {1{`RANDOM}};
  dataArray_58_4_cachedata_MPORT_en_pipe_0 = _RAND_2797[0:0];
  _RAND_2798 = {1{`RANDOM}};
  dataArray_58_4_cachedata_MPORT_addr_pipe_0 = _RAND_2798[1:0];
  _RAND_2800 = {1{`RANDOM}};
  dataArray_58_5_cachedata_MPORT_en_pipe_0 = _RAND_2800[0:0];
  _RAND_2801 = {1{`RANDOM}};
  dataArray_58_5_cachedata_MPORT_addr_pipe_0 = _RAND_2801[1:0];
  _RAND_2803 = {1{`RANDOM}};
  dataArray_58_6_cachedata_MPORT_en_pipe_0 = _RAND_2803[0:0];
  _RAND_2804 = {1{`RANDOM}};
  dataArray_58_6_cachedata_MPORT_addr_pipe_0 = _RAND_2804[1:0];
  _RAND_2806 = {1{`RANDOM}};
  dataArray_58_7_cachedata_MPORT_en_pipe_0 = _RAND_2806[0:0];
  _RAND_2807 = {1{`RANDOM}};
  dataArray_58_7_cachedata_MPORT_addr_pipe_0 = _RAND_2807[1:0];
  _RAND_2809 = {1{`RANDOM}};
  dataArray_58_8_cachedata_MPORT_en_pipe_0 = _RAND_2809[0:0];
  _RAND_2810 = {1{`RANDOM}};
  dataArray_58_8_cachedata_MPORT_addr_pipe_0 = _RAND_2810[1:0];
  _RAND_2812 = {1{`RANDOM}};
  dataArray_58_9_cachedata_MPORT_en_pipe_0 = _RAND_2812[0:0];
  _RAND_2813 = {1{`RANDOM}};
  dataArray_58_9_cachedata_MPORT_addr_pipe_0 = _RAND_2813[1:0];
  _RAND_2815 = {1{`RANDOM}};
  dataArray_58_10_cachedata_MPORT_en_pipe_0 = _RAND_2815[0:0];
  _RAND_2816 = {1{`RANDOM}};
  dataArray_58_10_cachedata_MPORT_addr_pipe_0 = _RAND_2816[1:0];
  _RAND_2818 = {1{`RANDOM}};
  dataArray_58_11_cachedata_MPORT_en_pipe_0 = _RAND_2818[0:0];
  _RAND_2819 = {1{`RANDOM}};
  dataArray_58_11_cachedata_MPORT_addr_pipe_0 = _RAND_2819[1:0];
  _RAND_2821 = {1{`RANDOM}};
  dataArray_58_12_cachedata_MPORT_en_pipe_0 = _RAND_2821[0:0];
  _RAND_2822 = {1{`RANDOM}};
  dataArray_58_12_cachedata_MPORT_addr_pipe_0 = _RAND_2822[1:0];
  _RAND_2824 = {1{`RANDOM}};
  dataArray_58_13_cachedata_MPORT_en_pipe_0 = _RAND_2824[0:0];
  _RAND_2825 = {1{`RANDOM}};
  dataArray_58_13_cachedata_MPORT_addr_pipe_0 = _RAND_2825[1:0];
  _RAND_2827 = {1{`RANDOM}};
  dataArray_58_14_cachedata_MPORT_en_pipe_0 = _RAND_2827[0:0];
  _RAND_2828 = {1{`RANDOM}};
  dataArray_58_14_cachedata_MPORT_addr_pipe_0 = _RAND_2828[1:0];
  _RAND_2830 = {1{`RANDOM}};
  dataArray_58_15_cachedata_MPORT_en_pipe_0 = _RAND_2830[0:0];
  _RAND_2831 = {1{`RANDOM}};
  dataArray_58_15_cachedata_MPORT_addr_pipe_0 = _RAND_2831[1:0];
  _RAND_2833 = {1{`RANDOM}};
  dataArray_59_0_cachedata_MPORT_en_pipe_0 = _RAND_2833[0:0];
  _RAND_2834 = {1{`RANDOM}};
  dataArray_59_0_cachedata_MPORT_addr_pipe_0 = _RAND_2834[1:0];
  _RAND_2836 = {1{`RANDOM}};
  dataArray_59_1_cachedata_MPORT_en_pipe_0 = _RAND_2836[0:0];
  _RAND_2837 = {1{`RANDOM}};
  dataArray_59_1_cachedata_MPORT_addr_pipe_0 = _RAND_2837[1:0];
  _RAND_2839 = {1{`RANDOM}};
  dataArray_59_2_cachedata_MPORT_en_pipe_0 = _RAND_2839[0:0];
  _RAND_2840 = {1{`RANDOM}};
  dataArray_59_2_cachedata_MPORT_addr_pipe_0 = _RAND_2840[1:0];
  _RAND_2842 = {1{`RANDOM}};
  dataArray_59_3_cachedata_MPORT_en_pipe_0 = _RAND_2842[0:0];
  _RAND_2843 = {1{`RANDOM}};
  dataArray_59_3_cachedata_MPORT_addr_pipe_0 = _RAND_2843[1:0];
  _RAND_2845 = {1{`RANDOM}};
  dataArray_59_4_cachedata_MPORT_en_pipe_0 = _RAND_2845[0:0];
  _RAND_2846 = {1{`RANDOM}};
  dataArray_59_4_cachedata_MPORT_addr_pipe_0 = _RAND_2846[1:0];
  _RAND_2848 = {1{`RANDOM}};
  dataArray_59_5_cachedata_MPORT_en_pipe_0 = _RAND_2848[0:0];
  _RAND_2849 = {1{`RANDOM}};
  dataArray_59_5_cachedata_MPORT_addr_pipe_0 = _RAND_2849[1:0];
  _RAND_2851 = {1{`RANDOM}};
  dataArray_59_6_cachedata_MPORT_en_pipe_0 = _RAND_2851[0:0];
  _RAND_2852 = {1{`RANDOM}};
  dataArray_59_6_cachedata_MPORT_addr_pipe_0 = _RAND_2852[1:0];
  _RAND_2854 = {1{`RANDOM}};
  dataArray_59_7_cachedata_MPORT_en_pipe_0 = _RAND_2854[0:0];
  _RAND_2855 = {1{`RANDOM}};
  dataArray_59_7_cachedata_MPORT_addr_pipe_0 = _RAND_2855[1:0];
  _RAND_2857 = {1{`RANDOM}};
  dataArray_59_8_cachedata_MPORT_en_pipe_0 = _RAND_2857[0:0];
  _RAND_2858 = {1{`RANDOM}};
  dataArray_59_8_cachedata_MPORT_addr_pipe_0 = _RAND_2858[1:0];
  _RAND_2860 = {1{`RANDOM}};
  dataArray_59_9_cachedata_MPORT_en_pipe_0 = _RAND_2860[0:0];
  _RAND_2861 = {1{`RANDOM}};
  dataArray_59_9_cachedata_MPORT_addr_pipe_0 = _RAND_2861[1:0];
  _RAND_2863 = {1{`RANDOM}};
  dataArray_59_10_cachedata_MPORT_en_pipe_0 = _RAND_2863[0:0];
  _RAND_2864 = {1{`RANDOM}};
  dataArray_59_10_cachedata_MPORT_addr_pipe_0 = _RAND_2864[1:0];
  _RAND_2866 = {1{`RANDOM}};
  dataArray_59_11_cachedata_MPORT_en_pipe_0 = _RAND_2866[0:0];
  _RAND_2867 = {1{`RANDOM}};
  dataArray_59_11_cachedata_MPORT_addr_pipe_0 = _RAND_2867[1:0];
  _RAND_2869 = {1{`RANDOM}};
  dataArray_59_12_cachedata_MPORT_en_pipe_0 = _RAND_2869[0:0];
  _RAND_2870 = {1{`RANDOM}};
  dataArray_59_12_cachedata_MPORT_addr_pipe_0 = _RAND_2870[1:0];
  _RAND_2872 = {1{`RANDOM}};
  dataArray_59_13_cachedata_MPORT_en_pipe_0 = _RAND_2872[0:0];
  _RAND_2873 = {1{`RANDOM}};
  dataArray_59_13_cachedata_MPORT_addr_pipe_0 = _RAND_2873[1:0];
  _RAND_2875 = {1{`RANDOM}};
  dataArray_59_14_cachedata_MPORT_en_pipe_0 = _RAND_2875[0:0];
  _RAND_2876 = {1{`RANDOM}};
  dataArray_59_14_cachedata_MPORT_addr_pipe_0 = _RAND_2876[1:0];
  _RAND_2878 = {1{`RANDOM}};
  dataArray_59_15_cachedata_MPORT_en_pipe_0 = _RAND_2878[0:0];
  _RAND_2879 = {1{`RANDOM}};
  dataArray_59_15_cachedata_MPORT_addr_pipe_0 = _RAND_2879[1:0];
  _RAND_2881 = {1{`RANDOM}};
  dataArray_60_0_cachedata_MPORT_en_pipe_0 = _RAND_2881[0:0];
  _RAND_2882 = {1{`RANDOM}};
  dataArray_60_0_cachedata_MPORT_addr_pipe_0 = _RAND_2882[1:0];
  _RAND_2884 = {1{`RANDOM}};
  dataArray_60_1_cachedata_MPORT_en_pipe_0 = _RAND_2884[0:0];
  _RAND_2885 = {1{`RANDOM}};
  dataArray_60_1_cachedata_MPORT_addr_pipe_0 = _RAND_2885[1:0];
  _RAND_2887 = {1{`RANDOM}};
  dataArray_60_2_cachedata_MPORT_en_pipe_0 = _RAND_2887[0:0];
  _RAND_2888 = {1{`RANDOM}};
  dataArray_60_2_cachedata_MPORT_addr_pipe_0 = _RAND_2888[1:0];
  _RAND_2890 = {1{`RANDOM}};
  dataArray_60_3_cachedata_MPORT_en_pipe_0 = _RAND_2890[0:0];
  _RAND_2891 = {1{`RANDOM}};
  dataArray_60_3_cachedata_MPORT_addr_pipe_0 = _RAND_2891[1:0];
  _RAND_2893 = {1{`RANDOM}};
  dataArray_60_4_cachedata_MPORT_en_pipe_0 = _RAND_2893[0:0];
  _RAND_2894 = {1{`RANDOM}};
  dataArray_60_4_cachedata_MPORT_addr_pipe_0 = _RAND_2894[1:0];
  _RAND_2896 = {1{`RANDOM}};
  dataArray_60_5_cachedata_MPORT_en_pipe_0 = _RAND_2896[0:0];
  _RAND_2897 = {1{`RANDOM}};
  dataArray_60_5_cachedata_MPORT_addr_pipe_0 = _RAND_2897[1:0];
  _RAND_2899 = {1{`RANDOM}};
  dataArray_60_6_cachedata_MPORT_en_pipe_0 = _RAND_2899[0:0];
  _RAND_2900 = {1{`RANDOM}};
  dataArray_60_6_cachedata_MPORT_addr_pipe_0 = _RAND_2900[1:0];
  _RAND_2902 = {1{`RANDOM}};
  dataArray_60_7_cachedata_MPORT_en_pipe_0 = _RAND_2902[0:0];
  _RAND_2903 = {1{`RANDOM}};
  dataArray_60_7_cachedata_MPORT_addr_pipe_0 = _RAND_2903[1:0];
  _RAND_2905 = {1{`RANDOM}};
  dataArray_60_8_cachedata_MPORT_en_pipe_0 = _RAND_2905[0:0];
  _RAND_2906 = {1{`RANDOM}};
  dataArray_60_8_cachedata_MPORT_addr_pipe_0 = _RAND_2906[1:0];
  _RAND_2908 = {1{`RANDOM}};
  dataArray_60_9_cachedata_MPORT_en_pipe_0 = _RAND_2908[0:0];
  _RAND_2909 = {1{`RANDOM}};
  dataArray_60_9_cachedata_MPORT_addr_pipe_0 = _RAND_2909[1:0];
  _RAND_2911 = {1{`RANDOM}};
  dataArray_60_10_cachedata_MPORT_en_pipe_0 = _RAND_2911[0:0];
  _RAND_2912 = {1{`RANDOM}};
  dataArray_60_10_cachedata_MPORT_addr_pipe_0 = _RAND_2912[1:0];
  _RAND_2914 = {1{`RANDOM}};
  dataArray_60_11_cachedata_MPORT_en_pipe_0 = _RAND_2914[0:0];
  _RAND_2915 = {1{`RANDOM}};
  dataArray_60_11_cachedata_MPORT_addr_pipe_0 = _RAND_2915[1:0];
  _RAND_2917 = {1{`RANDOM}};
  dataArray_60_12_cachedata_MPORT_en_pipe_0 = _RAND_2917[0:0];
  _RAND_2918 = {1{`RANDOM}};
  dataArray_60_12_cachedata_MPORT_addr_pipe_0 = _RAND_2918[1:0];
  _RAND_2920 = {1{`RANDOM}};
  dataArray_60_13_cachedata_MPORT_en_pipe_0 = _RAND_2920[0:0];
  _RAND_2921 = {1{`RANDOM}};
  dataArray_60_13_cachedata_MPORT_addr_pipe_0 = _RAND_2921[1:0];
  _RAND_2923 = {1{`RANDOM}};
  dataArray_60_14_cachedata_MPORT_en_pipe_0 = _RAND_2923[0:0];
  _RAND_2924 = {1{`RANDOM}};
  dataArray_60_14_cachedata_MPORT_addr_pipe_0 = _RAND_2924[1:0];
  _RAND_2926 = {1{`RANDOM}};
  dataArray_60_15_cachedata_MPORT_en_pipe_0 = _RAND_2926[0:0];
  _RAND_2927 = {1{`RANDOM}};
  dataArray_60_15_cachedata_MPORT_addr_pipe_0 = _RAND_2927[1:0];
  _RAND_2929 = {1{`RANDOM}};
  dataArray_61_0_cachedata_MPORT_en_pipe_0 = _RAND_2929[0:0];
  _RAND_2930 = {1{`RANDOM}};
  dataArray_61_0_cachedata_MPORT_addr_pipe_0 = _RAND_2930[1:0];
  _RAND_2932 = {1{`RANDOM}};
  dataArray_61_1_cachedata_MPORT_en_pipe_0 = _RAND_2932[0:0];
  _RAND_2933 = {1{`RANDOM}};
  dataArray_61_1_cachedata_MPORT_addr_pipe_0 = _RAND_2933[1:0];
  _RAND_2935 = {1{`RANDOM}};
  dataArray_61_2_cachedata_MPORT_en_pipe_0 = _RAND_2935[0:0];
  _RAND_2936 = {1{`RANDOM}};
  dataArray_61_2_cachedata_MPORT_addr_pipe_0 = _RAND_2936[1:0];
  _RAND_2938 = {1{`RANDOM}};
  dataArray_61_3_cachedata_MPORT_en_pipe_0 = _RAND_2938[0:0];
  _RAND_2939 = {1{`RANDOM}};
  dataArray_61_3_cachedata_MPORT_addr_pipe_0 = _RAND_2939[1:0];
  _RAND_2941 = {1{`RANDOM}};
  dataArray_61_4_cachedata_MPORT_en_pipe_0 = _RAND_2941[0:0];
  _RAND_2942 = {1{`RANDOM}};
  dataArray_61_4_cachedata_MPORT_addr_pipe_0 = _RAND_2942[1:0];
  _RAND_2944 = {1{`RANDOM}};
  dataArray_61_5_cachedata_MPORT_en_pipe_0 = _RAND_2944[0:0];
  _RAND_2945 = {1{`RANDOM}};
  dataArray_61_5_cachedata_MPORT_addr_pipe_0 = _RAND_2945[1:0];
  _RAND_2947 = {1{`RANDOM}};
  dataArray_61_6_cachedata_MPORT_en_pipe_0 = _RAND_2947[0:0];
  _RAND_2948 = {1{`RANDOM}};
  dataArray_61_6_cachedata_MPORT_addr_pipe_0 = _RAND_2948[1:0];
  _RAND_2950 = {1{`RANDOM}};
  dataArray_61_7_cachedata_MPORT_en_pipe_0 = _RAND_2950[0:0];
  _RAND_2951 = {1{`RANDOM}};
  dataArray_61_7_cachedata_MPORT_addr_pipe_0 = _RAND_2951[1:0];
  _RAND_2953 = {1{`RANDOM}};
  dataArray_61_8_cachedata_MPORT_en_pipe_0 = _RAND_2953[0:0];
  _RAND_2954 = {1{`RANDOM}};
  dataArray_61_8_cachedata_MPORT_addr_pipe_0 = _RAND_2954[1:0];
  _RAND_2956 = {1{`RANDOM}};
  dataArray_61_9_cachedata_MPORT_en_pipe_0 = _RAND_2956[0:0];
  _RAND_2957 = {1{`RANDOM}};
  dataArray_61_9_cachedata_MPORT_addr_pipe_0 = _RAND_2957[1:0];
  _RAND_2959 = {1{`RANDOM}};
  dataArray_61_10_cachedata_MPORT_en_pipe_0 = _RAND_2959[0:0];
  _RAND_2960 = {1{`RANDOM}};
  dataArray_61_10_cachedata_MPORT_addr_pipe_0 = _RAND_2960[1:0];
  _RAND_2962 = {1{`RANDOM}};
  dataArray_61_11_cachedata_MPORT_en_pipe_0 = _RAND_2962[0:0];
  _RAND_2963 = {1{`RANDOM}};
  dataArray_61_11_cachedata_MPORT_addr_pipe_0 = _RAND_2963[1:0];
  _RAND_2965 = {1{`RANDOM}};
  dataArray_61_12_cachedata_MPORT_en_pipe_0 = _RAND_2965[0:0];
  _RAND_2966 = {1{`RANDOM}};
  dataArray_61_12_cachedata_MPORT_addr_pipe_0 = _RAND_2966[1:0];
  _RAND_2968 = {1{`RANDOM}};
  dataArray_61_13_cachedata_MPORT_en_pipe_0 = _RAND_2968[0:0];
  _RAND_2969 = {1{`RANDOM}};
  dataArray_61_13_cachedata_MPORT_addr_pipe_0 = _RAND_2969[1:0];
  _RAND_2971 = {1{`RANDOM}};
  dataArray_61_14_cachedata_MPORT_en_pipe_0 = _RAND_2971[0:0];
  _RAND_2972 = {1{`RANDOM}};
  dataArray_61_14_cachedata_MPORT_addr_pipe_0 = _RAND_2972[1:0];
  _RAND_2974 = {1{`RANDOM}};
  dataArray_61_15_cachedata_MPORT_en_pipe_0 = _RAND_2974[0:0];
  _RAND_2975 = {1{`RANDOM}};
  dataArray_61_15_cachedata_MPORT_addr_pipe_0 = _RAND_2975[1:0];
  _RAND_2977 = {1{`RANDOM}};
  dataArray_62_0_cachedata_MPORT_en_pipe_0 = _RAND_2977[0:0];
  _RAND_2978 = {1{`RANDOM}};
  dataArray_62_0_cachedata_MPORT_addr_pipe_0 = _RAND_2978[1:0];
  _RAND_2980 = {1{`RANDOM}};
  dataArray_62_1_cachedata_MPORT_en_pipe_0 = _RAND_2980[0:0];
  _RAND_2981 = {1{`RANDOM}};
  dataArray_62_1_cachedata_MPORT_addr_pipe_0 = _RAND_2981[1:0];
  _RAND_2983 = {1{`RANDOM}};
  dataArray_62_2_cachedata_MPORT_en_pipe_0 = _RAND_2983[0:0];
  _RAND_2984 = {1{`RANDOM}};
  dataArray_62_2_cachedata_MPORT_addr_pipe_0 = _RAND_2984[1:0];
  _RAND_2986 = {1{`RANDOM}};
  dataArray_62_3_cachedata_MPORT_en_pipe_0 = _RAND_2986[0:0];
  _RAND_2987 = {1{`RANDOM}};
  dataArray_62_3_cachedata_MPORT_addr_pipe_0 = _RAND_2987[1:0];
  _RAND_2989 = {1{`RANDOM}};
  dataArray_62_4_cachedata_MPORT_en_pipe_0 = _RAND_2989[0:0];
  _RAND_2990 = {1{`RANDOM}};
  dataArray_62_4_cachedata_MPORT_addr_pipe_0 = _RAND_2990[1:0];
  _RAND_2992 = {1{`RANDOM}};
  dataArray_62_5_cachedata_MPORT_en_pipe_0 = _RAND_2992[0:0];
  _RAND_2993 = {1{`RANDOM}};
  dataArray_62_5_cachedata_MPORT_addr_pipe_0 = _RAND_2993[1:0];
  _RAND_2995 = {1{`RANDOM}};
  dataArray_62_6_cachedata_MPORT_en_pipe_0 = _RAND_2995[0:0];
  _RAND_2996 = {1{`RANDOM}};
  dataArray_62_6_cachedata_MPORT_addr_pipe_0 = _RAND_2996[1:0];
  _RAND_2998 = {1{`RANDOM}};
  dataArray_62_7_cachedata_MPORT_en_pipe_0 = _RAND_2998[0:0];
  _RAND_2999 = {1{`RANDOM}};
  dataArray_62_7_cachedata_MPORT_addr_pipe_0 = _RAND_2999[1:0];
  _RAND_3001 = {1{`RANDOM}};
  dataArray_62_8_cachedata_MPORT_en_pipe_0 = _RAND_3001[0:0];
  _RAND_3002 = {1{`RANDOM}};
  dataArray_62_8_cachedata_MPORT_addr_pipe_0 = _RAND_3002[1:0];
  _RAND_3004 = {1{`RANDOM}};
  dataArray_62_9_cachedata_MPORT_en_pipe_0 = _RAND_3004[0:0];
  _RAND_3005 = {1{`RANDOM}};
  dataArray_62_9_cachedata_MPORT_addr_pipe_0 = _RAND_3005[1:0];
  _RAND_3007 = {1{`RANDOM}};
  dataArray_62_10_cachedata_MPORT_en_pipe_0 = _RAND_3007[0:0];
  _RAND_3008 = {1{`RANDOM}};
  dataArray_62_10_cachedata_MPORT_addr_pipe_0 = _RAND_3008[1:0];
  _RAND_3010 = {1{`RANDOM}};
  dataArray_62_11_cachedata_MPORT_en_pipe_0 = _RAND_3010[0:0];
  _RAND_3011 = {1{`RANDOM}};
  dataArray_62_11_cachedata_MPORT_addr_pipe_0 = _RAND_3011[1:0];
  _RAND_3013 = {1{`RANDOM}};
  dataArray_62_12_cachedata_MPORT_en_pipe_0 = _RAND_3013[0:0];
  _RAND_3014 = {1{`RANDOM}};
  dataArray_62_12_cachedata_MPORT_addr_pipe_0 = _RAND_3014[1:0];
  _RAND_3016 = {1{`RANDOM}};
  dataArray_62_13_cachedata_MPORT_en_pipe_0 = _RAND_3016[0:0];
  _RAND_3017 = {1{`RANDOM}};
  dataArray_62_13_cachedata_MPORT_addr_pipe_0 = _RAND_3017[1:0];
  _RAND_3019 = {1{`RANDOM}};
  dataArray_62_14_cachedata_MPORT_en_pipe_0 = _RAND_3019[0:0];
  _RAND_3020 = {1{`RANDOM}};
  dataArray_62_14_cachedata_MPORT_addr_pipe_0 = _RAND_3020[1:0];
  _RAND_3022 = {1{`RANDOM}};
  dataArray_62_15_cachedata_MPORT_en_pipe_0 = _RAND_3022[0:0];
  _RAND_3023 = {1{`RANDOM}};
  dataArray_62_15_cachedata_MPORT_addr_pipe_0 = _RAND_3023[1:0];
  _RAND_3025 = {1{`RANDOM}};
  dataArray_63_0_cachedata_MPORT_en_pipe_0 = _RAND_3025[0:0];
  _RAND_3026 = {1{`RANDOM}};
  dataArray_63_0_cachedata_MPORT_addr_pipe_0 = _RAND_3026[1:0];
  _RAND_3028 = {1{`RANDOM}};
  dataArray_63_1_cachedata_MPORT_en_pipe_0 = _RAND_3028[0:0];
  _RAND_3029 = {1{`RANDOM}};
  dataArray_63_1_cachedata_MPORT_addr_pipe_0 = _RAND_3029[1:0];
  _RAND_3031 = {1{`RANDOM}};
  dataArray_63_2_cachedata_MPORT_en_pipe_0 = _RAND_3031[0:0];
  _RAND_3032 = {1{`RANDOM}};
  dataArray_63_2_cachedata_MPORT_addr_pipe_0 = _RAND_3032[1:0];
  _RAND_3034 = {1{`RANDOM}};
  dataArray_63_3_cachedata_MPORT_en_pipe_0 = _RAND_3034[0:0];
  _RAND_3035 = {1{`RANDOM}};
  dataArray_63_3_cachedata_MPORT_addr_pipe_0 = _RAND_3035[1:0];
  _RAND_3037 = {1{`RANDOM}};
  dataArray_63_4_cachedata_MPORT_en_pipe_0 = _RAND_3037[0:0];
  _RAND_3038 = {1{`RANDOM}};
  dataArray_63_4_cachedata_MPORT_addr_pipe_0 = _RAND_3038[1:0];
  _RAND_3040 = {1{`RANDOM}};
  dataArray_63_5_cachedata_MPORT_en_pipe_0 = _RAND_3040[0:0];
  _RAND_3041 = {1{`RANDOM}};
  dataArray_63_5_cachedata_MPORT_addr_pipe_0 = _RAND_3041[1:0];
  _RAND_3043 = {1{`RANDOM}};
  dataArray_63_6_cachedata_MPORT_en_pipe_0 = _RAND_3043[0:0];
  _RAND_3044 = {1{`RANDOM}};
  dataArray_63_6_cachedata_MPORT_addr_pipe_0 = _RAND_3044[1:0];
  _RAND_3046 = {1{`RANDOM}};
  dataArray_63_7_cachedata_MPORT_en_pipe_0 = _RAND_3046[0:0];
  _RAND_3047 = {1{`RANDOM}};
  dataArray_63_7_cachedata_MPORT_addr_pipe_0 = _RAND_3047[1:0];
  _RAND_3049 = {1{`RANDOM}};
  dataArray_63_8_cachedata_MPORT_en_pipe_0 = _RAND_3049[0:0];
  _RAND_3050 = {1{`RANDOM}};
  dataArray_63_8_cachedata_MPORT_addr_pipe_0 = _RAND_3050[1:0];
  _RAND_3052 = {1{`RANDOM}};
  dataArray_63_9_cachedata_MPORT_en_pipe_0 = _RAND_3052[0:0];
  _RAND_3053 = {1{`RANDOM}};
  dataArray_63_9_cachedata_MPORT_addr_pipe_0 = _RAND_3053[1:0];
  _RAND_3055 = {1{`RANDOM}};
  dataArray_63_10_cachedata_MPORT_en_pipe_0 = _RAND_3055[0:0];
  _RAND_3056 = {1{`RANDOM}};
  dataArray_63_10_cachedata_MPORT_addr_pipe_0 = _RAND_3056[1:0];
  _RAND_3058 = {1{`RANDOM}};
  dataArray_63_11_cachedata_MPORT_en_pipe_0 = _RAND_3058[0:0];
  _RAND_3059 = {1{`RANDOM}};
  dataArray_63_11_cachedata_MPORT_addr_pipe_0 = _RAND_3059[1:0];
  _RAND_3061 = {1{`RANDOM}};
  dataArray_63_12_cachedata_MPORT_en_pipe_0 = _RAND_3061[0:0];
  _RAND_3062 = {1{`RANDOM}};
  dataArray_63_12_cachedata_MPORT_addr_pipe_0 = _RAND_3062[1:0];
  _RAND_3064 = {1{`RANDOM}};
  dataArray_63_13_cachedata_MPORT_en_pipe_0 = _RAND_3064[0:0];
  _RAND_3065 = {1{`RANDOM}};
  dataArray_63_13_cachedata_MPORT_addr_pipe_0 = _RAND_3065[1:0];
  _RAND_3067 = {1{`RANDOM}};
  dataArray_63_14_cachedata_MPORT_en_pipe_0 = _RAND_3067[0:0];
  _RAND_3068 = {1{`RANDOM}};
  dataArray_63_14_cachedata_MPORT_addr_pipe_0 = _RAND_3068[1:0];
  _RAND_3070 = {1{`RANDOM}};
  dataArray_63_15_cachedata_MPORT_en_pipe_0 = _RAND_3070[0:0];
  _RAND_3071 = {1{`RANDOM}};
  dataArray_63_15_cachedata_MPORT_addr_pipe_0 = _RAND_3071[1:0];
  _RAND_3072 = {1{`RANDOM}};
  replace_set = _RAND_3072[1:0];
  _RAND_3073 = {1{`RANDOM}};
  random_num = _RAND_3073[1:0];
  _RAND_3074 = {1{`RANDOM}};
  tagArray_0_0 = _RAND_3074[19:0];
  _RAND_3075 = {1{`RANDOM}};
  tagArray_0_1 = _RAND_3075[19:0];
  _RAND_3076 = {1{`RANDOM}};
  tagArray_0_2 = _RAND_3076[19:0];
  _RAND_3077 = {1{`RANDOM}};
  tagArray_0_3 = _RAND_3077[19:0];
  _RAND_3078 = {1{`RANDOM}};
  tagArray_0_4 = _RAND_3078[19:0];
  _RAND_3079 = {1{`RANDOM}};
  tagArray_0_5 = _RAND_3079[19:0];
  _RAND_3080 = {1{`RANDOM}};
  tagArray_0_6 = _RAND_3080[19:0];
  _RAND_3081 = {1{`RANDOM}};
  tagArray_0_7 = _RAND_3081[19:0];
  _RAND_3082 = {1{`RANDOM}};
  tagArray_0_8 = _RAND_3082[19:0];
  _RAND_3083 = {1{`RANDOM}};
  tagArray_0_9 = _RAND_3083[19:0];
  _RAND_3084 = {1{`RANDOM}};
  tagArray_0_10 = _RAND_3084[19:0];
  _RAND_3085 = {1{`RANDOM}};
  tagArray_0_11 = _RAND_3085[19:0];
  _RAND_3086 = {1{`RANDOM}};
  tagArray_0_12 = _RAND_3086[19:0];
  _RAND_3087 = {1{`RANDOM}};
  tagArray_0_13 = _RAND_3087[19:0];
  _RAND_3088 = {1{`RANDOM}};
  tagArray_0_14 = _RAND_3088[19:0];
  _RAND_3089 = {1{`RANDOM}};
  tagArray_0_15 = _RAND_3089[19:0];
  _RAND_3090 = {1{`RANDOM}};
  tagArray_0_16 = _RAND_3090[19:0];
  _RAND_3091 = {1{`RANDOM}};
  tagArray_0_17 = _RAND_3091[19:0];
  _RAND_3092 = {1{`RANDOM}};
  tagArray_0_18 = _RAND_3092[19:0];
  _RAND_3093 = {1{`RANDOM}};
  tagArray_0_19 = _RAND_3093[19:0];
  _RAND_3094 = {1{`RANDOM}};
  tagArray_0_20 = _RAND_3094[19:0];
  _RAND_3095 = {1{`RANDOM}};
  tagArray_0_21 = _RAND_3095[19:0];
  _RAND_3096 = {1{`RANDOM}};
  tagArray_0_22 = _RAND_3096[19:0];
  _RAND_3097 = {1{`RANDOM}};
  tagArray_0_23 = _RAND_3097[19:0];
  _RAND_3098 = {1{`RANDOM}};
  tagArray_0_24 = _RAND_3098[19:0];
  _RAND_3099 = {1{`RANDOM}};
  tagArray_0_25 = _RAND_3099[19:0];
  _RAND_3100 = {1{`RANDOM}};
  tagArray_0_26 = _RAND_3100[19:0];
  _RAND_3101 = {1{`RANDOM}};
  tagArray_0_27 = _RAND_3101[19:0];
  _RAND_3102 = {1{`RANDOM}};
  tagArray_0_28 = _RAND_3102[19:0];
  _RAND_3103 = {1{`RANDOM}};
  tagArray_0_29 = _RAND_3103[19:0];
  _RAND_3104 = {1{`RANDOM}};
  tagArray_0_30 = _RAND_3104[19:0];
  _RAND_3105 = {1{`RANDOM}};
  tagArray_0_31 = _RAND_3105[19:0];
  _RAND_3106 = {1{`RANDOM}};
  tagArray_0_32 = _RAND_3106[19:0];
  _RAND_3107 = {1{`RANDOM}};
  tagArray_0_33 = _RAND_3107[19:0];
  _RAND_3108 = {1{`RANDOM}};
  tagArray_0_34 = _RAND_3108[19:0];
  _RAND_3109 = {1{`RANDOM}};
  tagArray_0_35 = _RAND_3109[19:0];
  _RAND_3110 = {1{`RANDOM}};
  tagArray_0_36 = _RAND_3110[19:0];
  _RAND_3111 = {1{`RANDOM}};
  tagArray_0_37 = _RAND_3111[19:0];
  _RAND_3112 = {1{`RANDOM}};
  tagArray_0_38 = _RAND_3112[19:0];
  _RAND_3113 = {1{`RANDOM}};
  tagArray_0_39 = _RAND_3113[19:0];
  _RAND_3114 = {1{`RANDOM}};
  tagArray_0_40 = _RAND_3114[19:0];
  _RAND_3115 = {1{`RANDOM}};
  tagArray_0_41 = _RAND_3115[19:0];
  _RAND_3116 = {1{`RANDOM}};
  tagArray_0_42 = _RAND_3116[19:0];
  _RAND_3117 = {1{`RANDOM}};
  tagArray_0_43 = _RAND_3117[19:0];
  _RAND_3118 = {1{`RANDOM}};
  tagArray_0_44 = _RAND_3118[19:0];
  _RAND_3119 = {1{`RANDOM}};
  tagArray_0_45 = _RAND_3119[19:0];
  _RAND_3120 = {1{`RANDOM}};
  tagArray_0_46 = _RAND_3120[19:0];
  _RAND_3121 = {1{`RANDOM}};
  tagArray_0_47 = _RAND_3121[19:0];
  _RAND_3122 = {1{`RANDOM}};
  tagArray_0_48 = _RAND_3122[19:0];
  _RAND_3123 = {1{`RANDOM}};
  tagArray_0_49 = _RAND_3123[19:0];
  _RAND_3124 = {1{`RANDOM}};
  tagArray_0_50 = _RAND_3124[19:0];
  _RAND_3125 = {1{`RANDOM}};
  tagArray_0_51 = _RAND_3125[19:0];
  _RAND_3126 = {1{`RANDOM}};
  tagArray_0_52 = _RAND_3126[19:0];
  _RAND_3127 = {1{`RANDOM}};
  tagArray_0_53 = _RAND_3127[19:0];
  _RAND_3128 = {1{`RANDOM}};
  tagArray_0_54 = _RAND_3128[19:0];
  _RAND_3129 = {1{`RANDOM}};
  tagArray_0_55 = _RAND_3129[19:0];
  _RAND_3130 = {1{`RANDOM}};
  tagArray_0_56 = _RAND_3130[19:0];
  _RAND_3131 = {1{`RANDOM}};
  tagArray_0_57 = _RAND_3131[19:0];
  _RAND_3132 = {1{`RANDOM}};
  tagArray_0_58 = _RAND_3132[19:0];
  _RAND_3133 = {1{`RANDOM}};
  tagArray_0_59 = _RAND_3133[19:0];
  _RAND_3134 = {1{`RANDOM}};
  tagArray_0_60 = _RAND_3134[19:0];
  _RAND_3135 = {1{`RANDOM}};
  tagArray_0_61 = _RAND_3135[19:0];
  _RAND_3136 = {1{`RANDOM}};
  tagArray_0_62 = _RAND_3136[19:0];
  _RAND_3137 = {1{`RANDOM}};
  tagArray_0_63 = _RAND_3137[19:0];
  _RAND_3138 = {1{`RANDOM}};
  tagArray_1_0 = _RAND_3138[19:0];
  _RAND_3139 = {1{`RANDOM}};
  tagArray_1_1 = _RAND_3139[19:0];
  _RAND_3140 = {1{`RANDOM}};
  tagArray_1_2 = _RAND_3140[19:0];
  _RAND_3141 = {1{`RANDOM}};
  tagArray_1_3 = _RAND_3141[19:0];
  _RAND_3142 = {1{`RANDOM}};
  tagArray_1_4 = _RAND_3142[19:0];
  _RAND_3143 = {1{`RANDOM}};
  tagArray_1_5 = _RAND_3143[19:0];
  _RAND_3144 = {1{`RANDOM}};
  tagArray_1_6 = _RAND_3144[19:0];
  _RAND_3145 = {1{`RANDOM}};
  tagArray_1_7 = _RAND_3145[19:0];
  _RAND_3146 = {1{`RANDOM}};
  tagArray_1_8 = _RAND_3146[19:0];
  _RAND_3147 = {1{`RANDOM}};
  tagArray_1_9 = _RAND_3147[19:0];
  _RAND_3148 = {1{`RANDOM}};
  tagArray_1_10 = _RAND_3148[19:0];
  _RAND_3149 = {1{`RANDOM}};
  tagArray_1_11 = _RAND_3149[19:0];
  _RAND_3150 = {1{`RANDOM}};
  tagArray_1_12 = _RAND_3150[19:0];
  _RAND_3151 = {1{`RANDOM}};
  tagArray_1_13 = _RAND_3151[19:0];
  _RAND_3152 = {1{`RANDOM}};
  tagArray_1_14 = _RAND_3152[19:0];
  _RAND_3153 = {1{`RANDOM}};
  tagArray_1_15 = _RAND_3153[19:0];
  _RAND_3154 = {1{`RANDOM}};
  tagArray_1_16 = _RAND_3154[19:0];
  _RAND_3155 = {1{`RANDOM}};
  tagArray_1_17 = _RAND_3155[19:0];
  _RAND_3156 = {1{`RANDOM}};
  tagArray_1_18 = _RAND_3156[19:0];
  _RAND_3157 = {1{`RANDOM}};
  tagArray_1_19 = _RAND_3157[19:0];
  _RAND_3158 = {1{`RANDOM}};
  tagArray_1_20 = _RAND_3158[19:0];
  _RAND_3159 = {1{`RANDOM}};
  tagArray_1_21 = _RAND_3159[19:0];
  _RAND_3160 = {1{`RANDOM}};
  tagArray_1_22 = _RAND_3160[19:0];
  _RAND_3161 = {1{`RANDOM}};
  tagArray_1_23 = _RAND_3161[19:0];
  _RAND_3162 = {1{`RANDOM}};
  tagArray_1_24 = _RAND_3162[19:0];
  _RAND_3163 = {1{`RANDOM}};
  tagArray_1_25 = _RAND_3163[19:0];
  _RAND_3164 = {1{`RANDOM}};
  tagArray_1_26 = _RAND_3164[19:0];
  _RAND_3165 = {1{`RANDOM}};
  tagArray_1_27 = _RAND_3165[19:0];
  _RAND_3166 = {1{`RANDOM}};
  tagArray_1_28 = _RAND_3166[19:0];
  _RAND_3167 = {1{`RANDOM}};
  tagArray_1_29 = _RAND_3167[19:0];
  _RAND_3168 = {1{`RANDOM}};
  tagArray_1_30 = _RAND_3168[19:0];
  _RAND_3169 = {1{`RANDOM}};
  tagArray_1_31 = _RAND_3169[19:0];
  _RAND_3170 = {1{`RANDOM}};
  tagArray_1_32 = _RAND_3170[19:0];
  _RAND_3171 = {1{`RANDOM}};
  tagArray_1_33 = _RAND_3171[19:0];
  _RAND_3172 = {1{`RANDOM}};
  tagArray_1_34 = _RAND_3172[19:0];
  _RAND_3173 = {1{`RANDOM}};
  tagArray_1_35 = _RAND_3173[19:0];
  _RAND_3174 = {1{`RANDOM}};
  tagArray_1_36 = _RAND_3174[19:0];
  _RAND_3175 = {1{`RANDOM}};
  tagArray_1_37 = _RAND_3175[19:0];
  _RAND_3176 = {1{`RANDOM}};
  tagArray_1_38 = _RAND_3176[19:0];
  _RAND_3177 = {1{`RANDOM}};
  tagArray_1_39 = _RAND_3177[19:0];
  _RAND_3178 = {1{`RANDOM}};
  tagArray_1_40 = _RAND_3178[19:0];
  _RAND_3179 = {1{`RANDOM}};
  tagArray_1_41 = _RAND_3179[19:0];
  _RAND_3180 = {1{`RANDOM}};
  tagArray_1_42 = _RAND_3180[19:0];
  _RAND_3181 = {1{`RANDOM}};
  tagArray_1_43 = _RAND_3181[19:0];
  _RAND_3182 = {1{`RANDOM}};
  tagArray_1_44 = _RAND_3182[19:0];
  _RAND_3183 = {1{`RANDOM}};
  tagArray_1_45 = _RAND_3183[19:0];
  _RAND_3184 = {1{`RANDOM}};
  tagArray_1_46 = _RAND_3184[19:0];
  _RAND_3185 = {1{`RANDOM}};
  tagArray_1_47 = _RAND_3185[19:0];
  _RAND_3186 = {1{`RANDOM}};
  tagArray_1_48 = _RAND_3186[19:0];
  _RAND_3187 = {1{`RANDOM}};
  tagArray_1_49 = _RAND_3187[19:0];
  _RAND_3188 = {1{`RANDOM}};
  tagArray_1_50 = _RAND_3188[19:0];
  _RAND_3189 = {1{`RANDOM}};
  tagArray_1_51 = _RAND_3189[19:0];
  _RAND_3190 = {1{`RANDOM}};
  tagArray_1_52 = _RAND_3190[19:0];
  _RAND_3191 = {1{`RANDOM}};
  tagArray_1_53 = _RAND_3191[19:0];
  _RAND_3192 = {1{`RANDOM}};
  tagArray_1_54 = _RAND_3192[19:0];
  _RAND_3193 = {1{`RANDOM}};
  tagArray_1_55 = _RAND_3193[19:0];
  _RAND_3194 = {1{`RANDOM}};
  tagArray_1_56 = _RAND_3194[19:0];
  _RAND_3195 = {1{`RANDOM}};
  tagArray_1_57 = _RAND_3195[19:0];
  _RAND_3196 = {1{`RANDOM}};
  tagArray_1_58 = _RAND_3196[19:0];
  _RAND_3197 = {1{`RANDOM}};
  tagArray_1_59 = _RAND_3197[19:0];
  _RAND_3198 = {1{`RANDOM}};
  tagArray_1_60 = _RAND_3198[19:0];
  _RAND_3199 = {1{`RANDOM}};
  tagArray_1_61 = _RAND_3199[19:0];
  _RAND_3200 = {1{`RANDOM}};
  tagArray_1_62 = _RAND_3200[19:0];
  _RAND_3201 = {1{`RANDOM}};
  tagArray_1_63 = _RAND_3201[19:0];
  _RAND_3202 = {1{`RANDOM}};
  tagArray_2_0 = _RAND_3202[19:0];
  _RAND_3203 = {1{`RANDOM}};
  tagArray_2_1 = _RAND_3203[19:0];
  _RAND_3204 = {1{`RANDOM}};
  tagArray_2_2 = _RAND_3204[19:0];
  _RAND_3205 = {1{`RANDOM}};
  tagArray_2_3 = _RAND_3205[19:0];
  _RAND_3206 = {1{`RANDOM}};
  tagArray_2_4 = _RAND_3206[19:0];
  _RAND_3207 = {1{`RANDOM}};
  tagArray_2_5 = _RAND_3207[19:0];
  _RAND_3208 = {1{`RANDOM}};
  tagArray_2_6 = _RAND_3208[19:0];
  _RAND_3209 = {1{`RANDOM}};
  tagArray_2_7 = _RAND_3209[19:0];
  _RAND_3210 = {1{`RANDOM}};
  tagArray_2_8 = _RAND_3210[19:0];
  _RAND_3211 = {1{`RANDOM}};
  tagArray_2_9 = _RAND_3211[19:0];
  _RAND_3212 = {1{`RANDOM}};
  tagArray_2_10 = _RAND_3212[19:0];
  _RAND_3213 = {1{`RANDOM}};
  tagArray_2_11 = _RAND_3213[19:0];
  _RAND_3214 = {1{`RANDOM}};
  tagArray_2_12 = _RAND_3214[19:0];
  _RAND_3215 = {1{`RANDOM}};
  tagArray_2_13 = _RAND_3215[19:0];
  _RAND_3216 = {1{`RANDOM}};
  tagArray_2_14 = _RAND_3216[19:0];
  _RAND_3217 = {1{`RANDOM}};
  tagArray_2_15 = _RAND_3217[19:0];
  _RAND_3218 = {1{`RANDOM}};
  tagArray_2_16 = _RAND_3218[19:0];
  _RAND_3219 = {1{`RANDOM}};
  tagArray_2_17 = _RAND_3219[19:0];
  _RAND_3220 = {1{`RANDOM}};
  tagArray_2_18 = _RAND_3220[19:0];
  _RAND_3221 = {1{`RANDOM}};
  tagArray_2_19 = _RAND_3221[19:0];
  _RAND_3222 = {1{`RANDOM}};
  tagArray_2_20 = _RAND_3222[19:0];
  _RAND_3223 = {1{`RANDOM}};
  tagArray_2_21 = _RAND_3223[19:0];
  _RAND_3224 = {1{`RANDOM}};
  tagArray_2_22 = _RAND_3224[19:0];
  _RAND_3225 = {1{`RANDOM}};
  tagArray_2_23 = _RAND_3225[19:0];
  _RAND_3226 = {1{`RANDOM}};
  tagArray_2_24 = _RAND_3226[19:0];
  _RAND_3227 = {1{`RANDOM}};
  tagArray_2_25 = _RAND_3227[19:0];
  _RAND_3228 = {1{`RANDOM}};
  tagArray_2_26 = _RAND_3228[19:0];
  _RAND_3229 = {1{`RANDOM}};
  tagArray_2_27 = _RAND_3229[19:0];
  _RAND_3230 = {1{`RANDOM}};
  tagArray_2_28 = _RAND_3230[19:0];
  _RAND_3231 = {1{`RANDOM}};
  tagArray_2_29 = _RAND_3231[19:0];
  _RAND_3232 = {1{`RANDOM}};
  tagArray_2_30 = _RAND_3232[19:0];
  _RAND_3233 = {1{`RANDOM}};
  tagArray_2_31 = _RAND_3233[19:0];
  _RAND_3234 = {1{`RANDOM}};
  tagArray_2_32 = _RAND_3234[19:0];
  _RAND_3235 = {1{`RANDOM}};
  tagArray_2_33 = _RAND_3235[19:0];
  _RAND_3236 = {1{`RANDOM}};
  tagArray_2_34 = _RAND_3236[19:0];
  _RAND_3237 = {1{`RANDOM}};
  tagArray_2_35 = _RAND_3237[19:0];
  _RAND_3238 = {1{`RANDOM}};
  tagArray_2_36 = _RAND_3238[19:0];
  _RAND_3239 = {1{`RANDOM}};
  tagArray_2_37 = _RAND_3239[19:0];
  _RAND_3240 = {1{`RANDOM}};
  tagArray_2_38 = _RAND_3240[19:0];
  _RAND_3241 = {1{`RANDOM}};
  tagArray_2_39 = _RAND_3241[19:0];
  _RAND_3242 = {1{`RANDOM}};
  tagArray_2_40 = _RAND_3242[19:0];
  _RAND_3243 = {1{`RANDOM}};
  tagArray_2_41 = _RAND_3243[19:0];
  _RAND_3244 = {1{`RANDOM}};
  tagArray_2_42 = _RAND_3244[19:0];
  _RAND_3245 = {1{`RANDOM}};
  tagArray_2_43 = _RAND_3245[19:0];
  _RAND_3246 = {1{`RANDOM}};
  tagArray_2_44 = _RAND_3246[19:0];
  _RAND_3247 = {1{`RANDOM}};
  tagArray_2_45 = _RAND_3247[19:0];
  _RAND_3248 = {1{`RANDOM}};
  tagArray_2_46 = _RAND_3248[19:0];
  _RAND_3249 = {1{`RANDOM}};
  tagArray_2_47 = _RAND_3249[19:0];
  _RAND_3250 = {1{`RANDOM}};
  tagArray_2_48 = _RAND_3250[19:0];
  _RAND_3251 = {1{`RANDOM}};
  tagArray_2_49 = _RAND_3251[19:0];
  _RAND_3252 = {1{`RANDOM}};
  tagArray_2_50 = _RAND_3252[19:0];
  _RAND_3253 = {1{`RANDOM}};
  tagArray_2_51 = _RAND_3253[19:0];
  _RAND_3254 = {1{`RANDOM}};
  tagArray_2_52 = _RAND_3254[19:0];
  _RAND_3255 = {1{`RANDOM}};
  tagArray_2_53 = _RAND_3255[19:0];
  _RAND_3256 = {1{`RANDOM}};
  tagArray_2_54 = _RAND_3256[19:0];
  _RAND_3257 = {1{`RANDOM}};
  tagArray_2_55 = _RAND_3257[19:0];
  _RAND_3258 = {1{`RANDOM}};
  tagArray_2_56 = _RAND_3258[19:0];
  _RAND_3259 = {1{`RANDOM}};
  tagArray_2_57 = _RAND_3259[19:0];
  _RAND_3260 = {1{`RANDOM}};
  tagArray_2_58 = _RAND_3260[19:0];
  _RAND_3261 = {1{`RANDOM}};
  tagArray_2_59 = _RAND_3261[19:0];
  _RAND_3262 = {1{`RANDOM}};
  tagArray_2_60 = _RAND_3262[19:0];
  _RAND_3263 = {1{`RANDOM}};
  tagArray_2_61 = _RAND_3263[19:0];
  _RAND_3264 = {1{`RANDOM}};
  tagArray_2_62 = _RAND_3264[19:0];
  _RAND_3265 = {1{`RANDOM}};
  tagArray_2_63 = _RAND_3265[19:0];
  _RAND_3266 = {1{`RANDOM}};
  tagArray_3_0 = _RAND_3266[19:0];
  _RAND_3267 = {1{`RANDOM}};
  tagArray_3_1 = _RAND_3267[19:0];
  _RAND_3268 = {1{`RANDOM}};
  tagArray_3_2 = _RAND_3268[19:0];
  _RAND_3269 = {1{`RANDOM}};
  tagArray_3_3 = _RAND_3269[19:0];
  _RAND_3270 = {1{`RANDOM}};
  tagArray_3_4 = _RAND_3270[19:0];
  _RAND_3271 = {1{`RANDOM}};
  tagArray_3_5 = _RAND_3271[19:0];
  _RAND_3272 = {1{`RANDOM}};
  tagArray_3_6 = _RAND_3272[19:0];
  _RAND_3273 = {1{`RANDOM}};
  tagArray_3_7 = _RAND_3273[19:0];
  _RAND_3274 = {1{`RANDOM}};
  tagArray_3_8 = _RAND_3274[19:0];
  _RAND_3275 = {1{`RANDOM}};
  tagArray_3_9 = _RAND_3275[19:0];
  _RAND_3276 = {1{`RANDOM}};
  tagArray_3_10 = _RAND_3276[19:0];
  _RAND_3277 = {1{`RANDOM}};
  tagArray_3_11 = _RAND_3277[19:0];
  _RAND_3278 = {1{`RANDOM}};
  tagArray_3_12 = _RAND_3278[19:0];
  _RAND_3279 = {1{`RANDOM}};
  tagArray_3_13 = _RAND_3279[19:0];
  _RAND_3280 = {1{`RANDOM}};
  tagArray_3_14 = _RAND_3280[19:0];
  _RAND_3281 = {1{`RANDOM}};
  tagArray_3_15 = _RAND_3281[19:0];
  _RAND_3282 = {1{`RANDOM}};
  tagArray_3_16 = _RAND_3282[19:0];
  _RAND_3283 = {1{`RANDOM}};
  tagArray_3_17 = _RAND_3283[19:0];
  _RAND_3284 = {1{`RANDOM}};
  tagArray_3_18 = _RAND_3284[19:0];
  _RAND_3285 = {1{`RANDOM}};
  tagArray_3_19 = _RAND_3285[19:0];
  _RAND_3286 = {1{`RANDOM}};
  tagArray_3_20 = _RAND_3286[19:0];
  _RAND_3287 = {1{`RANDOM}};
  tagArray_3_21 = _RAND_3287[19:0];
  _RAND_3288 = {1{`RANDOM}};
  tagArray_3_22 = _RAND_3288[19:0];
  _RAND_3289 = {1{`RANDOM}};
  tagArray_3_23 = _RAND_3289[19:0];
  _RAND_3290 = {1{`RANDOM}};
  tagArray_3_24 = _RAND_3290[19:0];
  _RAND_3291 = {1{`RANDOM}};
  tagArray_3_25 = _RAND_3291[19:0];
  _RAND_3292 = {1{`RANDOM}};
  tagArray_3_26 = _RAND_3292[19:0];
  _RAND_3293 = {1{`RANDOM}};
  tagArray_3_27 = _RAND_3293[19:0];
  _RAND_3294 = {1{`RANDOM}};
  tagArray_3_28 = _RAND_3294[19:0];
  _RAND_3295 = {1{`RANDOM}};
  tagArray_3_29 = _RAND_3295[19:0];
  _RAND_3296 = {1{`RANDOM}};
  tagArray_3_30 = _RAND_3296[19:0];
  _RAND_3297 = {1{`RANDOM}};
  tagArray_3_31 = _RAND_3297[19:0];
  _RAND_3298 = {1{`RANDOM}};
  tagArray_3_32 = _RAND_3298[19:0];
  _RAND_3299 = {1{`RANDOM}};
  tagArray_3_33 = _RAND_3299[19:0];
  _RAND_3300 = {1{`RANDOM}};
  tagArray_3_34 = _RAND_3300[19:0];
  _RAND_3301 = {1{`RANDOM}};
  tagArray_3_35 = _RAND_3301[19:0];
  _RAND_3302 = {1{`RANDOM}};
  tagArray_3_36 = _RAND_3302[19:0];
  _RAND_3303 = {1{`RANDOM}};
  tagArray_3_37 = _RAND_3303[19:0];
  _RAND_3304 = {1{`RANDOM}};
  tagArray_3_38 = _RAND_3304[19:0];
  _RAND_3305 = {1{`RANDOM}};
  tagArray_3_39 = _RAND_3305[19:0];
  _RAND_3306 = {1{`RANDOM}};
  tagArray_3_40 = _RAND_3306[19:0];
  _RAND_3307 = {1{`RANDOM}};
  tagArray_3_41 = _RAND_3307[19:0];
  _RAND_3308 = {1{`RANDOM}};
  tagArray_3_42 = _RAND_3308[19:0];
  _RAND_3309 = {1{`RANDOM}};
  tagArray_3_43 = _RAND_3309[19:0];
  _RAND_3310 = {1{`RANDOM}};
  tagArray_3_44 = _RAND_3310[19:0];
  _RAND_3311 = {1{`RANDOM}};
  tagArray_3_45 = _RAND_3311[19:0];
  _RAND_3312 = {1{`RANDOM}};
  tagArray_3_46 = _RAND_3312[19:0];
  _RAND_3313 = {1{`RANDOM}};
  tagArray_3_47 = _RAND_3313[19:0];
  _RAND_3314 = {1{`RANDOM}};
  tagArray_3_48 = _RAND_3314[19:0];
  _RAND_3315 = {1{`RANDOM}};
  tagArray_3_49 = _RAND_3315[19:0];
  _RAND_3316 = {1{`RANDOM}};
  tagArray_3_50 = _RAND_3316[19:0];
  _RAND_3317 = {1{`RANDOM}};
  tagArray_3_51 = _RAND_3317[19:0];
  _RAND_3318 = {1{`RANDOM}};
  tagArray_3_52 = _RAND_3318[19:0];
  _RAND_3319 = {1{`RANDOM}};
  tagArray_3_53 = _RAND_3319[19:0];
  _RAND_3320 = {1{`RANDOM}};
  tagArray_3_54 = _RAND_3320[19:0];
  _RAND_3321 = {1{`RANDOM}};
  tagArray_3_55 = _RAND_3321[19:0];
  _RAND_3322 = {1{`RANDOM}};
  tagArray_3_56 = _RAND_3322[19:0];
  _RAND_3323 = {1{`RANDOM}};
  tagArray_3_57 = _RAND_3323[19:0];
  _RAND_3324 = {1{`RANDOM}};
  tagArray_3_58 = _RAND_3324[19:0];
  _RAND_3325 = {1{`RANDOM}};
  tagArray_3_59 = _RAND_3325[19:0];
  _RAND_3326 = {1{`RANDOM}};
  tagArray_3_60 = _RAND_3326[19:0];
  _RAND_3327 = {1{`RANDOM}};
  tagArray_3_61 = _RAND_3327[19:0];
  _RAND_3328 = {1{`RANDOM}};
  tagArray_3_62 = _RAND_3328[19:0];
  _RAND_3329 = {1{`RANDOM}};
  tagArray_3_63 = _RAND_3329[19:0];
  _RAND_3330 = {1{`RANDOM}};
  validArray_0_0 = _RAND_3330[0:0];
  _RAND_3331 = {1{`RANDOM}};
  validArray_0_1 = _RAND_3331[0:0];
  _RAND_3332 = {1{`RANDOM}};
  validArray_0_2 = _RAND_3332[0:0];
  _RAND_3333 = {1{`RANDOM}};
  validArray_0_3 = _RAND_3333[0:0];
  _RAND_3334 = {1{`RANDOM}};
  validArray_0_4 = _RAND_3334[0:0];
  _RAND_3335 = {1{`RANDOM}};
  validArray_0_5 = _RAND_3335[0:0];
  _RAND_3336 = {1{`RANDOM}};
  validArray_0_6 = _RAND_3336[0:0];
  _RAND_3337 = {1{`RANDOM}};
  validArray_0_7 = _RAND_3337[0:0];
  _RAND_3338 = {1{`RANDOM}};
  validArray_0_8 = _RAND_3338[0:0];
  _RAND_3339 = {1{`RANDOM}};
  validArray_0_9 = _RAND_3339[0:0];
  _RAND_3340 = {1{`RANDOM}};
  validArray_0_10 = _RAND_3340[0:0];
  _RAND_3341 = {1{`RANDOM}};
  validArray_0_11 = _RAND_3341[0:0];
  _RAND_3342 = {1{`RANDOM}};
  validArray_0_12 = _RAND_3342[0:0];
  _RAND_3343 = {1{`RANDOM}};
  validArray_0_13 = _RAND_3343[0:0];
  _RAND_3344 = {1{`RANDOM}};
  validArray_0_14 = _RAND_3344[0:0];
  _RAND_3345 = {1{`RANDOM}};
  validArray_0_15 = _RAND_3345[0:0];
  _RAND_3346 = {1{`RANDOM}};
  validArray_0_16 = _RAND_3346[0:0];
  _RAND_3347 = {1{`RANDOM}};
  validArray_0_17 = _RAND_3347[0:0];
  _RAND_3348 = {1{`RANDOM}};
  validArray_0_18 = _RAND_3348[0:0];
  _RAND_3349 = {1{`RANDOM}};
  validArray_0_19 = _RAND_3349[0:0];
  _RAND_3350 = {1{`RANDOM}};
  validArray_0_20 = _RAND_3350[0:0];
  _RAND_3351 = {1{`RANDOM}};
  validArray_0_21 = _RAND_3351[0:0];
  _RAND_3352 = {1{`RANDOM}};
  validArray_0_22 = _RAND_3352[0:0];
  _RAND_3353 = {1{`RANDOM}};
  validArray_0_23 = _RAND_3353[0:0];
  _RAND_3354 = {1{`RANDOM}};
  validArray_0_24 = _RAND_3354[0:0];
  _RAND_3355 = {1{`RANDOM}};
  validArray_0_25 = _RAND_3355[0:0];
  _RAND_3356 = {1{`RANDOM}};
  validArray_0_26 = _RAND_3356[0:0];
  _RAND_3357 = {1{`RANDOM}};
  validArray_0_27 = _RAND_3357[0:0];
  _RAND_3358 = {1{`RANDOM}};
  validArray_0_28 = _RAND_3358[0:0];
  _RAND_3359 = {1{`RANDOM}};
  validArray_0_29 = _RAND_3359[0:0];
  _RAND_3360 = {1{`RANDOM}};
  validArray_0_30 = _RAND_3360[0:0];
  _RAND_3361 = {1{`RANDOM}};
  validArray_0_31 = _RAND_3361[0:0];
  _RAND_3362 = {1{`RANDOM}};
  validArray_0_32 = _RAND_3362[0:0];
  _RAND_3363 = {1{`RANDOM}};
  validArray_0_33 = _RAND_3363[0:0];
  _RAND_3364 = {1{`RANDOM}};
  validArray_0_34 = _RAND_3364[0:0];
  _RAND_3365 = {1{`RANDOM}};
  validArray_0_35 = _RAND_3365[0:0];
  _RAND_3366 = {1{`RANDOM}};
  validArray_0_36 = _RAND_3366[0:0];
  _RAND_3367 = {1{`RANDOM}};
  validArray_0_37 = _RAND_3367[0:0];
  _RAND_3368 = {1{`RANDOM}};
  validArray_0_38 = _RAND_3368[0:0];
  _RAND_3369 = {1{`RANDOM}};
  validArray_0_39 = _RAND_3369[0:0];
  _RAND_3370 = {1{`RANDOM}};
  validArray_0_40 = _RAND_3370[0:0];
  _RAND_3371 = {1{`RANDOM}};
  validArray_0_41 = _RAND_3371[0:0];
  _RAND_3372 = {1{`RANDOM}};
  validArray_0_42 = _RAND_3372[0:0];
  _RAND_3373 = {1{`RANDOM}};
  validArray_0_43 = _RAND_3373[0:0];
  _RAND_3374 = {1{`RANDOM}};
  validArray_0_44 = _RAND_3374[0:0];
  _RAND_3375 = {1{`RANDOM}};
  validArray_0_45 = _RAND_3375[0:0];
  _RAND_3376 = {1{`RANDOM}};
  validArray_0_46 = _RAND_3376[0:0];
  _RAND_3377 = {1{`RANDOM}};
  validArray_0_47 = _RAND_3377[0:0];
  _RAND_3378 = {1{`RANDOM}};
  validArray_0_48 = _RAND_3378[0:0];
  _RAND_3379 = {1{`RANDOM}};
  validArray_0_49 = _RAND_3379[0:0];
  _RAND_3380 = {1{`RANDOM}};
  validArray_0_50 = _RAND_3380[0:0];
  _RAND_3381 = {1{`RANDOM}};
  validArray_0_51 = _RAND_3381[0:0];
  _RAND_3382 = {1{`RANDOM}};
  validArray_0_52 = _RAND_3382[0:0];
  _RAND_3383 = {1{`RANDOM}};
  validArray_0_53 = _RAND_3383[0:0];
  _RAND_3384 = {1{`RANDOM}};
  validArray_0_54 = _RAND_3384[0:0];
  _RAND_3385 = {1{`RANDOM}};
  validArray_0_55 = _RAND_3385[0:0];
  _RAND_3386 = {1{`RANDOM}};
  validArray_0_56 = _RAND_3386[0:0];
  _RAND_3387 = {1{`RANDOM}};
  validArray_0_57 = _RAND_3387[0:0];
  _RAND_3388 = {1{`RANDOM}};
  validArray_0_58 = _RAND_3388[0:0];
  _RAND_3389 = {1{`RANDOM}};
  validArray_0_59 = _RAND_3389[0:0];
  _RAND_3390 = {1{`RANDOM}};
  validArray_0_60 = _RAND_3390[0:0];
  _RAND_3391 = {1{`RANDOM}};
  validArray_0_61 = _RAND_3391[0:0];
  _RAND_3392 = {1{`RANDOM}};
  validArray_0_62 = _RAND_3392[0:0];
  _RAND_3393 = {1{`RANDOM}};
  validArray_0_63 = _RAND_3393[0:0];
  _RAND_3394 = {1{`RANDOM}};
  validArray_1_0 = _RAND_3394[0:0];
  _RAND_3395 = {1{`RANDOM}};
  validArray_1_1 = _RAND_3395[0:0];
  _RAND_3396 = {1{`RANDOM}};
  validArray_1_2 = _RAND_3396[0:0];
  _RAND_3397 = {1{`RANDOM}};
  validArray_1_3 = _RAND_3397[0:0];
  _RAND_3398 = {1{`RANDOM}};
  validArray_1_4 = _RAND_3398[0:0];
  _RAND_3399 = {1{`RANDOM}};
  validArray_1_5 = _RAND_3399[0:0];
  _RAND_3400 = {1{`RANDOM}};
  validArray_1_6 = _RAND_3400[0:0];
  _RAND_3401 = {1{`RANDOM}};
  validArray_1_7 = _RAND_3401[0:0];
  _RAND_3402 = {1{`RANDOM}};
  validArray_1_8 = _RAND_3402[0:0];
  _RAND_3403 = {1{`RANDOM}};
  validArray_1_9 = _RAND_3403[0:0];
  _RAND_3404 = {1{`RANDOM}};
  validArray_1_10 = _RAND_3404[0:0];
  _RAND_3405 = {1{`RANDOM}};
  validArray_1_11 = _RAND_3405[0:0];
  _RAND_3406 = {1{`RANDOM}};
  validArray_1_12 = _RAND_3406[0:0];
  _RAND_3407 = {1{`RANDOM}};
  validArray_1_13 = _RAND_3407[0:0];
  _RAND_3408 = {1{`RANDOM}};
  validArray_1_14 = _RAND_3408[0:0];
  _RAND_3409 = {1{`RANDOM}};
  validArray_1_15 = _RAND_3409[0:0];
  _RAND_3410 = {1{`RANDOM}};
  validArray_1_16 = _RAND_3410[0:0];
  _RAND_3411 = {1{`RANDOM}};
  validArray_1_17 = _RAND_3411[0:0];
  _RAND_3412 = {1{`RANDOM}};
  validArray_1_18 = _RAND_3412[0:0];
  _RAND_3413 = {1{`RANDOM}};
  validArray_1_19 = _RAND_3413[0:0];
  _RAND_3414 = {1{`RANDOM}};
  validArray_1_20 = _RAND_3414[0:0];
  _RAND_3415 = {1{`RANDOM}};
  validArray_1_21 = _RAND_3415[0:0];
  _RAND_3416 = {1{`RANDOM}};
  validArray_1_22 = _RAND_3416[0:0];
  _RAND_3417 = {1{`RANDOM}};
  validArray_1_23 = _RAND_3417[0:0];
  _RAND_3418 = {1{`RANDOM}};
  validArray_1_24 = _RAND_3418[0:0];
  _RAND_3419 = {1{`RANDOM}};
  validArray_1_25 = _RAND_3419[0:0];
  _RAND_3420 = {1{`RANDOM}};
  validArray_1_26 = _RAND_3420[0:0];
  _RAND_3421 = {1{`RANDOM}};
  validArray_1_27 = _RAND_3421[0:0];
  _RAND_3422 = {1{`RANDOM}};
  validArray_1_28 = _RAND_3422[0:0];
  _RAND_3423 = {1{`RANDOM}};
  validArray_1_29 = _RAND_3423[0:0];
  _RAND_3424 = {1{`RANDOM}};
  validArray_1_30 = _RAND_3424[0:0];
  _RAND_3425 = {1{`RANDOM}};
  validArray_1_31 = _RAND_3425[0:0];
  _RAND_3426 = {1{`RANDOM}};
  validArray_1_32 = _RAND_3426[0:0];
  _RAND_3427 = {1{`RANDOM}};
  validArray_1_33 = _RAND_3427[0:0];
  _RAND_3428 = {1{`RANDOM}};
  validArray_1_34 = _RAND_3428[0:0];
  _RAND_3429 = {1{`RANDOM}};
  validArray_1_35 = _RAND_3429[0:0];
  _RAND_3430 = {1{`RANDOM}};
  validArray_1_36 = _RAND_3430[0:0];
  _RAND_3431 = {1{`RANDOM}};
  validArray_1_37 = _RAND_3431[0:0];
  _RAND_3432 = {1{`RANDOM}};
  validArray_1_38 = _RAND_3432[0:0];
  _RAND_3433 = {1{`RANDOM}};
  validArray_1_39 = _RAND_3433[0:0];
  _RAND_3434 = {1{`RANDOM}};
  validArray_1_40 = _RAND_3434[0:0];
  _RAND_3435 = {1{`RANDOM}};
  validArray_1_41 = _RAND_3435[0:0];
  _RAND_3436 = {1{`RANDOM}};
  validArray_1_42 = _RAND_3436[0:0];
  _RAND_3437 = {1{`RANDOM}};
  validArray_1_43 = _RAND_3437[0:0];
  _RAND_3438 = {1{`RANDOM}};
  validArray_1_44 = _RAND_3438[0:0];
  _RAND_3439 = {1{`RANDOM}};
  validArray_1_45 = _RAND_3439[0:0];
  _RAND_3440 = {1{`RANDOM}};
  validArray_1_46 = _RAND_3440[0:0];
  _RAND_3441 = {1{`RANDOM}};
  validArray_1_47 = _RAND_3441[0:0];
  _RAND_3442 = {1{`RANDOM}};
  validArray_1_48 = _RAND_3442[0:0];
  _RAND_3443 = {1{`RANDOM}};
  validArray_1_49 = _RAND_3443[0:0];
  _RAND_3444 = {1{`RANDOM}};
  validArray_1_50 = _RAND_3444[0:0];
  _RAND_3445 = {1{`RANDOM}};
  validArray_1_51 = _RAND_3445[0:0];
  _RAND_3446 = {1{`RANDOM}};
  validArray_1_52 = _RAND_3446[0:0];
  _RAND_3447 = {1{`RANDOM}};
  validArray_1_53 = _RAND_3447[0:0];
  _RAND_3448 = {1{`RANDOM}};
  validArray_1_54 = _RAND_3448[0:0];
  _RAND_3449 = {1{`RANDOM}};
  validArray_1_55 = _RAND_3449[0:0];
  _RAND_3450 = {1{`RANDOM}};
  validArray_1_56 = _RAND_3450[0:0];
  _RAND_3451 = {1{`RANDOM}};
  validArray_1_57 = _RAND_3451[0:0];
  _RAND_3452 = {1{`RANDOM}};
  validArray_1_58 = _RAND_3452[0:0];
  _RAND_3453 = {1{`RANDOM}};
  validArray_1_59 = _RAND_3453[0:0];
  _RAND_3454 = {1{`RANDOM}};
  validArray_1_60 = _RAND_3454[0:0];
  _RAND_3455 = {1{`RANDOM}};
  validArray_1_61 = _RAND_3455[0:0];
  _RAND_3456 = {1{`RANDOM}};
  validArray_1_62 = _RAND_3456[0:0];
  _RAND_3457 = {1{`RANDOM}};
  validArray_1_63 = _RAND_3457[0:0];
  _RAND_3458 = {1{`RANDOM}};
  validArray_2_0 = _RAND_3458[0:0];
  _RAND_3459 = {1{`RANDOM}};
  validArray_2_1 = _RAND_3459[0:0];
  _RAND_3460 = {1{`RANDOM}};
  validArray_2_2 = _RAND_3460[0:0];
  _RAND_3461 = {1{`RANDOM}};
  validArray_2_3 = _RAND_3461[0:0];
  _RAND_3462 = {1{`RANDOM}};
  validArray_2_4 = _RAND_3462[0:0];
  _RAND_3463 = {1{`RANDOM}};
  validArray_2_5 = _RAND_3463[0:0];
  _RAND_3464 = {1{`RANDOM}};
  validArray_2_6 = _RAND_3464[0:0];
  _RAND_3465 = {1{`RANDOM}};
  validArray_2_7 = _RAND_3465[0:0];
  _RAND_3466 = {1{`RANDOM}};
  validArray_2_8 = _RAND_3466[0:0];
  _RAND_3467 = {1{`RANDOM}};
  validArray_2_9 = _RAND_3467[0:0];
  _RAND_3468 = {1{`RANDOM}};
  validArray_2_10 = _RAND_3468[0:0];
  _RAND_3469 = {1{`RANDOM}};
  validArray_2_11 = _RAND_3469[0:0];
  _RAND_3470 = {1{`RANDOM}};
  validArray_2_12 = _RAND_3470[0:0];
  _RAND_3471 = {1{`RANDOM}};
  validArray_2_13 = _RAND_3471[0:0];
  _RAND_3472 = {1{`RANDOM}};
  validArray_2_14 = _RAND_3472[0:0];
  _RAND_3473 = {1{`RANDOM}};
  validArray_2_15 = _RAND_3473[0:0];
  _RAND_3474 = {1{`RANDOM}};
  validArray_2_16 = _RAND_3474[0:0];
  _RAND_3475 = {1{`RANDOM}};
  validArray_2_17 = _RAND_3475[0:0];
  _RAND_3476 = {1{`RANDOM}};
  validArray_2_18 = _RAND_3476[0:0];
  _RAND_3477 = {1{`RANDOM}};
  validArray_2_19 = _RAND_3477[0:0];
  _RAND_3478 = {1{`RANDOM}};
  validArray_2_20 = _RAND_3478[0:0];
  _RAND_3479 = {1{`RANDOM}};
  validArray_2_21 = _RAND_3479[0:0];
  _RAND_3480 = {1{`RANDOM}};
  validArray_2_22 = _RAND_3480[0:0];
  _RAND_3481 = {1{`RANDOM}};
  validArray_2_23 = _RAND_3481[0:0];
  _RAND_3482 = {1{`RANDOM}};
  validArray_2_24 = _RAND_3482[0:0];
  _RAND_3483 = {1{`RANDOM}};
  validArray_2_25 = _RAND_3483[0:0];
  _RAND_3484 = {1{`RANDOM}};
  validArray_2_26 = _RAND_3484[0:0];
  _RAND_3485 = {1{`RANDOM}};
  validArray_2_27 = _RAND_3485[0:0];
  _RAND_3486 = {1{`RANDOM}};
  validArray_2_28 = _RAND_3486[0:0];
  _RAND_3487 = {1{`RANDOM}};
  validArray_2_29 = _RAND_3487[0:0];
  _RAND_3488 = {1{`RANDOM}};
  validArray_2_30 = _RAND_3488[0:0];
  _RAND_3489 = {1{`RANDOM}};
  validArray_2_31 = _RAND_3489[0:0];
  _RAND_3490 = {1{`RANDOM}};
  validArray_2_32 = _RAND_3490[0:0];
  _RAND_3491 = {1{`RANDOM}};
  validArray_2_33 = _RAND_3491[0:0];
  _RAND_3492 = {1{`RANDOM}};
  validArray_2_34 = _RAND_3492[0:0];
  _RAND_3493 = {1{`RANDOM}};
  validArray_2_35 = _RAND_3493[0:0];
  _RAND_3494 = {1{`RANDOM}};
  validArray_2_36 = _RAND_3494[0:0];
  _RAND_3495 = {1{`RANDOM}};
  validArray_2_37 = _RAND_3495[0:0];
  _RAND_3496 = {1{`RANDOM}};
  validArray_2_38 = _RAND_3496[0:0];
  _RAND_3497 = {1{`RANDOM}};
  validArray_2_39 = _RAND_3497[0:0];
  _RAND_3498 = {1{`RANDOM}};
  validArray_2_40 = _RAND_3498[0:0];
  _RAND_3499 = {1{`RANDOM}};
  validArray_2_41 = _RAND_3499[0:0];
  _RAND_3500 = {1{`RANDOM}};
  validArray_2_42 = _RAND_3500[0:0];
  _RAND_3501 = {1{`RANDOM}};
  validArray_2_43 = _RAND_3501[0:0];
  _RAND_3502 = {1{`RANDOM}};
  validArray_2_44 = _RAND_3502[0:0];
  _RAND_3503 = {1{`RANDOM}};
  validArray_2_45 = _RAND_3503[0:0];
  _RAND_3504 = {1{`RANDOM}};
  validArray_2_46 = _RAND_3504[0:0];
  _RAND_3505 = {1{`RANDOM}};
  validArray_2_47 = _RAND_3505[0:0];
  _RAND_3506 = {1{`RANDOM}};
  validArray_2_48 = _RAND_3506[0:0];
  _RAND_3507 = {1{`RANDOM}};
  validArray_2_49 = _RAND_3507[0:0];
  _RAND_3508 = {1{`RANDOM}};
  validArray_2_50 = _RAND_3508[0:0];
  _RAND_3509 = {1{`RANDOM}};
  validArray_2_51 = _RAND_3509[0:0];
  _RAND_3510 = {1{`RANDOM}};
  validArray_2_52 = _RAND_3510[0:0];
  _RAND_3511 = {1{`RANDOM}};
  validArray_2_53 = _RAND_3511[0:0];
  _RAND_3512 = {1{`RANDOM}};
  validArray_2_54 = _RAND_3512[0:0];
  _RAND_3513 = {1{`RANDOM}};
  validArray_2_55 = _RAND_3513[0:0];
  _RAND_3514 = {1{`RANDOM}};
  validArray_2_56 = _RAND_3514[0:0];
  _RAND_3515 = {1{`RANDOM}};
  validArray_2_57 = _RAND_3515[0:0];
  _RAND_3516 = {1{`RANDOM}};
  validArray_2_58 = _RAND_3516[0:0];
  _RAND_3517 = {1{`RANDOM}};
  validArray_2_59 = _RAND_3517[0:0];
  _RAND_3518 = {1{`RANDOM}};
  validArray_2_60 = _RAND_3518[0:0];
  _RAND_3519 = {1{`RANDOM}};
  validArray_2_61 = _RAND_3519[0:0];
  _RAND_3520 = {1{`RANDOM}};
  validArray_2_62 = _RAND_3520[0:0];
  _RAND_3521 = {1{`RANDOM}};
  validArray_2_63 = _RAND_3521[0:0];
  _RAND_3522 = {1{`RANDOM}};
  validArray_3_0 = _RAND_3522[0:0];
  _RAND_3523 = {1{`RANDOM}};
  validArray_3_1 = _RAND_3523[0:0];
  _RAND_3524 = {1{`RANDOM}};
  validArray_3_2 = _RAND_3524[0:0];
  _RAND_3525 = {1{`RANDOM}};
  validArray_3_3 = _RAND_3525[0:0];
  _RAND_3526 = {1{`RANDOM}};
  validArray_3_4 = _RAND_3526[0:0];
  _RAND_3527 = {1{`RANDOM}};
  validArray_3_5 = _RAND_3527[0:0];
  _RAND_3528 = {1{`RANDOM}};
  validArray_3_6 = _RAND_3528[0:0];
  _RAND_3529 = {1{`RANDOM}};
  validArray_3_7 = _RAND_3529[0:0];
  _RAND_3530 = {1{`RANDOM}};
  validArray_3_8 = _RAND_3530[0:0];
  _RAND_3531 = {1{`RANDOM}};
  validArray_3_9 = _RAND_3531[0:0];
  _RAND_3532 = {1{`RANDOM}};
  validArray_3_10 = _RAND_3532[0:0];
  _RAND_3533 = {1{`RANDOM}};
  validArray_3_11 = _RAND_3533[0:0];
  _RAND_3534 = {1{`RANDOM}};
  validArray_3_12 = _RAND_3534[0:0];
  _RAND_3535 = {1{`RANDOM}};
  validArray_3_13 = _RAND_3535[0:0];
  _RAND_3536 = {1{`RANDOM}};
  validArray_3_14 = _RAND_3536[0:0];
  _RAND_3537 = {1{`RANDOM}};
  validArray_3_15 = _RAND_3537[0:0];
  _RAND_3538 = {1{`RANDOM}};
  validArray_3_16 = _RAND_3538[0:0];
  _RAND_3539 = {1{`RANDOM}};
  validArray_3_17 = _RAND_3539[0:0];
  _RAND_3540 = {1{`RANDOM}};
  validArray_3_18 = _RAND_3540[0:0];
  _RAND_3541 = {1{`RANDOM}};
  validArray_3_19 = _RAND_3541[0:0];
  _RAND_3542 = {1{`RANDOM}};
  validArray_3_20 = _RAND_3542[0:0];
  _RAND_3543 = {1{`RANDOM}};
  validArray_3_21 = _RAND_3543[0:0];
  _RAND_3544 = {1{`RANDOM}};
  validArray_3_22 = _RAND_3544[0:0];
  _RAND_3545 = {1{`RANDOM}};
  validArray_3_23 = _RAND_3545[0:0];
  _RAND_3546 = {1{`RANDOM}};
  validArray_3_24 = _RAND_3546[0:0];
  _RAND_3547 = {1{`RANDOM}};
  validArray_3_25 = _RAND_3547[0:0];
  _RAND_3548 = {1{`RANDOM}};
  validArray_3_26 = _RAND_3548[0:0];
  _RAND_3549 = {1{`RANDOM}};
  validArray_3_27 = _RAND_3549[0:0];
  _RAND_3550 = {1{`RANDOM}};
  validArray_3_28 = _RAND_3550[0:0];
  _RAND_3551 = {1{`RANDOM}};
  validArray_3_29 = _RAND_3551[0:0];
  _RAND_3552 = {1{`RANDOM}};
  validArray_3_30 = _RAND_3552[0:0];
  _RAND_3553 = {1{`RANDOM}};
  validArray_3_31 = _RAND_3553[0:0];
  _RAND_3554 = {1{`RANDOM}};
  validArray_3_32 = _RAND_3554[0:0];
  _RAND_3555 = {1{`RANDOM}};
  validArray_3_33 = _RAND_3555[0:0];
  _RAND_3556 = {1{`RANDOM}};
  validArray_3_34 = _RAND_3556[0:0];
  _RAND_3557 = {1{`RANDOM}};
  validArray_3_35 = _RAND_3557[0:0];
  _RAND_3558 = {1{`RANDOM}};
  validArray_3_36 = _RAND_3558[0:0];
  _RAND_3559 = {1{`RANDOM}};
  validArray_3_37 = _RAND_3559[0:0];
  _RAND_3560 = {1{`RANDOM}};
  validArray_3_38 = _RAND_3560[0:0];
  _RAND_3561 = {1{`RANDOM}};
  validArray_3_39 = _RAND_3561[0:0];
  _RAND_3562 = {1{`RANDOM}};
  validArray_3_40 = _RAND_3562[0:0];
  _RAND_3563 = {1{`RANDOM}};
  validArray_3_41 = _RAND_3563[0:0];
  _RAND_3564 = {1{`RANDOM}};
  validArray_3_42 = _RAND_3564[0:0];
  _RAND_3565 = {1{`RANDOM}};
  validArray_3_43 = _RAND_3565[0:0];
  _RAND_3566 = {1{`RANDOM}};
  validArray_3_44 = _RAND_3566[0:0];
  _RAND_3567 = {1{`RANDOM}};
  validArray_3_45 = _RAND_3567[0:0];
  _RAND_3568 = {1{`RANDOM}};
  validArray_3_46 = _RAND_3568[0:0];
  _RAND_3569 = {1{`RANDOM}};
  validArray_3_47 = _RAND_3569[0:0];
  _RAND_3570 = {1{`RANDOM}};
  validArray_3_48 = _RAND_3570[0:0];
  _RAND_3571 = {1{`RANDOM}};
  validArray_3_49 = _RAND_3571[0:0];
  _RAND_3572 = {1{`RANDOM}};
  validArray_3_50 = _RAND_3572[0:0];
  _RAND_3573 = {1{`RANDOM}};
  validArray_3_51 = _RAND_3573[0:0];
  _RAND_3574 = {1{`RANDOM}};
  validArray_3_52 = _RAND_3574[0:0];
  _RAND_3575 = {1{`RANDOM}};
  validArray_3_53 = _RAND_3575[0:0];
  _RAND_3576 = {1{`RANDOM}};
  validArray_3_54 = _RAND_3576[0:0];
  _RAND_3577 = {1{`RANDOM}};
  validArray_3_55 = _RAND_3577[0:0];
  _RAND_3578 = {1{`RANDOM}};
  validArray_3_56 = _RAND_3578[0:0];
  _RAND_3579 = {1{`RANDOM}};
  validArray_3_57 = _RAND_3579[0:0];
  _RAND_3580 = {1{`RANDOM}};
  validArray_3_58 = _RAND_3580[0:0];
  _RAND_3581 = {1{`RANDOM}};
  validArray_3_59 = _RAND_3581[0:0];
  _RAND_3582 = {1{`RANDOM}};
  validArray_3_60 = _RAND_3582[0:0];
  _RAND_3583 = {1{`RANDOM}};
  validArray_3_61 = _RAND_3583[0:0];
  _RAND_3584 = {1{`RANDOM}};
  validArray_3_62 = _RAND_3584[0:0];
  _RAND_3585 = {1{`RANDOM}};
  validArray_3_63 = _RAND_3585[0:0];
  _RAND_3586 = {1{`RANDOM}};
  off = _RAND_3586[3:0];
  _RAND_3587 = {1{`RANDOM}};
  state_cache = _RAND_3587[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAM_axi(
  input         clock,
  input         reset,
  output        axi_ar_ready,
  input         axi_ar_valid,
  input  [31:0] axi_ar_bits_addr,
  input  [7:0]  axi_ar_bits_len,
  input         axi_r_ready,
  output        axi_r_valid,
  output [31:0] axi_r_bits_data,
  output        axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  RamBB_i1_clock; // @[sram_Axi.scala 65:26]
  wire [31:0] RamBB_i1_addr; // @[sram_Axi.scala 65:26]
  wire  RamBB_i1_mem_wen; // @[sram_Axi.scala 65:26]
  wire  RamBB_i1_valid; // @[sram_Axi.scala 65:26]
  wire [31:0] RamBB_i1_wdata; // @[sram_Axi.scala 65:26]
  wire [3:0] RamBB_i1_wmask; // @[sram_Axi.scala 65:26]
  wire [31:0] RamBB_i1_rdata; // @[sram_Axi.scala 65:26]
  reg  delay; // @[sram_Axi.scala 22:24]
  reg [7:0] reg_AxLen; // @[sram_Axi.scala 25:28]
  reg [31:0] reg_addr; // @[sram_Axi.scala 26:28]
  reg [1:0] reg_burst; // @[sram_Axi.scala 27:28]
  reg [1:0] state_sram; // @[sram_Axi.scala 31:29]
  wire  _T_1 = axi_ar_ready & axi_ar_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_sram_T_1 = reg_AxLen == 8'h0 ? 2'h3 : 2'h2; // @[sram_Axi.scala 47:34]
  wire  _T_4 = 2'h2 == state_sram; // @[sram_Axi.scala 32:25]
  wire [1:0] _state_sram_T_3 = reg_AxLen == 8'h1 ? 2'h3 : 2'h2; // @[sram_Axi.scala 54:31]
  wire  _reg_AxLen_T = axi_r_ready & axi_r_valid; // @[Decoupled.scala 51:35]
  wire [7:0] _reg_AxLen_T_2 = reg_AxLen - 8'h1; // @[sram_Axi.scala 55:53]
  wire [7:0] _reg_AxLen_T_3 = _reg_AxLen_T ? _reg_AxLen_T_2 : reg_AxLen; // @[sram_Axi.scala 55:31]
  wire [31:0] _reg_addr_T_2 = reg_addr + 32'h4; // @[sram_Axi.scala 57:53]
  wire [31:0] _reg_addr_T_3 = _reg_AxLen_T ? _reg_addr_T_2 : reg_addr; // @[sram_Axi.scala 57:30]
  wire [31:0] _reg_addr_T_5 = 2'h1 == reg_burst ? _reg_addr_T_3 : reg_addr; // @[Mux.scala 81:58]
  wire  _T_5 = 2'h3 == state_sram; // @[sram_Axi.scala 32:25]
  wire [1:0] _GEN_5 = 2'h3 == state_sram ? 2'h0 : state_sram; // @[sram_Axi.scala 32:25 61:24 31:29]
  RamBB RamBB_i1 ( // @[sram_Axi.scala 65:26]
    .clock(RamBB_i1_clock),
    .addr(RamBB_i1_addr),
    .mem_wen(RamBB_i1_mem_wen),
    .valid(RamBB_i1_valid),
    .wdata(RamBB_i1_wdata),
    .wmask(RamBB_i1_wmask),
    .rdata(RamBB_i1_rdata)
  );
  assign axi_ar_ready = 2'h0 == state_sram; // @[Mux.scala 81:61]
  assign axi_r_valid = _T_5 | _T_4; // @[Mux.scala 81:58]
  assign axi_r_bits_data = RamBB_i1_rdata; // @[sram_Axi.scala 78:21]
  assign axi_r_bits_last = state_sram == 2'h3; // @[sram_Axi.scala 80:39]
  assign RamBB_i1_clock = clock; // @[sram_Axi.scala 66:25]
  assign RamBB_i1_addr = reg_addr; // @[sram_Axi.scala 67:25]
  assign RamBB_i1_mem_wen = 1'h0; // @[sram_Axi.scala 68:25]
  assign RamBB_i1_valid = _T_5 | _T_4; // @[Mux.scala 81:58]
  assign RamBB_i1_wdata = 32'h0; // @[sram_Axi.scala 72:25]
  assign RamBB_i1_wmask = 4'h0; // @[sram_Axi.scala 73:25]
  always @(posedge clock) begin
    if (reset) begin // @[sram_Axi.scala 22:24]
      delay <= 1'h0; // @[sram_Axi.scala 22:24]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      delay <= 1'h0; // @[sram_Axi.scala 34:19]
    end else if (2'h1 == state_sram) begin // @[sram_Axi.scala 32:25]
      delay <= delay - 1'h1; // @[sram_Axi.scala 51:19]
    end
    if (reset) begin // @[sram_Axi.scala 25:28]
      reg_AxLen <= 8'h0; // @[sram_Axi.scala 25:28]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        reg_AxLen <= axi_ar_bits_len; // @[sram_Axi.scala 38:28]
      end
    end else if (!(2'h1 == state_sram)) begin // @[sram_Axi.scala 32:25]
      if (2'h2 == state_sram) begin // @[sram_Axi.scala 32:25]
        reg_AxLen <= _reg_AxLen_T_3; // @[sram_Axi.scala 55:25]
      end
    end
    if (reset) begin // @[sram_Axi.scala 26:28]
      reg_addr <= 32'h0; // @[sram_Axi.scala 26:28]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        reg_addr <= axi_ar_bits_addr; // @[sram_Axi.scala 39:28]
      end
    end else if (!(2'h1 == state_sram)) begin // @[sram_Axi.scala 32:25]
      if (2'h2 == state_sram) begin // @[sram_Axi.scala 32:25]
        reg_addr <= _reg_addr_T_5; // @[sram_Axi.scala 56:25]
      end
    end
    if (reset) begin // @[sram_Axi.scala 27:28]
      reg_burst <= 2'h3; // @[sram_Axi.scala 27:28]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        reg_burst <= 2'h1; // @[sram_Axi.scala 40:28]
      end
    end
    if (reset) begin // @[sram_Axi.scala 31:29]
      state_sram <= 2'h0; // @[sram_Axi.scala 31:29]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        state_sram <= 2'h1; // @[sram_Axi.scala 37:28]
      end else begin
        state_sram <= 2'h0; // @[sram_Axi.scala 42:28]
      end
    end else if (2'h1 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (~delay) begin // @[sram_Axi.scala 46:34]
        state_sram <= _state_sram_T_1; // @[sram_Axi.scala 47:28]
      end else begin
        state_sram <= 2'h1; // @[sram_Axi.scala 49:28]
      end
    end else if (2'h2 == state_sram) begin // @[sram_Axi.scala 32:25]
      state_sram <= _state_sram_T_3; // @[sram_Axi.scala 54:25]
    end else begin
      state_sram <= _GEN_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_AxLen = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  reg_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_burst = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  state_sram = _RAND_4[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAM(
  input         clock,
  input         reset,
  output        axi_ar_ready,
  input         axi_ar_valid,
  input  [31:0] axi_ar_bits_addr,
  input         axi_r_ready,
  output        axi_r_valid,
  output [31:0] axi_r_bits_data,
  output        axi_aw_ready,
  input         axi_aw_valid,
  input  [31:0] axi_aw_bits_addr,
  output        axi_w_ready,
  input         axi_w_valid,
  input  [31:0] axi_w_bits_data,
  input  [3:0]  axi_w_bits_strb,
  input         axi_b_ready,
  output        axi_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RamBB_i1_clock; // @[sram_AxiLite.scala 77:26]
  wire [31:0] RamBB_i1_addr; // @[sram_AxiLite.scala 77:26]
  wire  RamBB_i1_mem_wen; // @[sram_AxiLite.scala 77:26]
  wire  RamBB_i1_valid; // @[sram_AxiLite.scala 77:26]
  wire [31:0] RamBB_i1_wdata; // @[sram_AxiLite.scala 77:26]
  wire [3:0] RamBB_i1_wmask; // @[sram_AxiLite.scala 77:26]
  wire [31:0] RamBB_i1_rdata; // @[sram_AxiLite.scala 77:26]
  reg  delay; // @[sram_AxiLite.scala 42:24]
  reg [2:0] state; // @[sram_AxiLite.scala 46:24]
  wire  _T_1 = axi_ar_ready & axi_ar_valid; // @[Decoupled.scala 51:35]
  wire  _T_2 = axi_aw_ready & axi_aw_valid; // @[Decoupled.scala 51:35]
  wire  _T_3 = axi_w_ready & axi_w_valid; // @[Decoupled.scala 51:35]
  wire  _state_T = ~delay; // @[sram_AxiLite.scala 62:32]
  wire  _delay_T_1 = delay - 1'h1; // @[sram_AxiLite.scala 63:28]
  wire  _T_6 = 3'h2 == state; // @[sram_AxiLite.scala 47:20]
  wire  _state_T_2 = axi_r_ready & axi_r_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_3 = _state_T_2 ? 3'h0 : 3'h2; // @[sram_AxiLite.scala 66:25]
  wire [2:0] _state_T_5 = _state_T ? 3'h4 : 3'h3; // @[sram_AxiLite.scala 69:25]
  wire  _T_8 = 3'h4 == state; // @[sram_AxiLite.scala 47:20]
  wire  _state_T_6 = axi_b_ready & axi_b_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_7 = _state_T_6 ? 3'h0 : 3'h4; // @[sram_AxiLite.scala 73:25]
  wire [2:0] _GEN_2 = 3'h4 == state ? _state_T_7 : state; // @[sram_AxiLite.scala 47:20 73:19 46:24]
  wire [2:0] _GEN_3 = 3'h3 == state ? _state_T_5 : _GEN_2; // @[sram_AxiLite.scala 47:20 69:19]
  wire  _GEN_4 = 3'h3 == state ? _delay_T_1 : delay; // @[sram_AxiLite.scala 47:20 70:19 42:24]
  wire [31:0] _RamBB_i1_io_addr_T_1 = _T_6 ? axi_ar_bits_addr : 32'h0; // @[Mux.scala 81:58]
  RamBB RamBB_i1 ( // @[sram_AxiLite.scala 77:26]
    .clock(RamBB_i1_clock),
    .addr(RamBB_i1_addr),
    .mem_wen(RamBB_i1_mem_wen),
    .valid(RamBB_i1_valid),
    .wdata(RamBB_i1_wdata),
    .wmask(RamBB_i1_wmask),
    .rdata(RamBB_i1_rdata)
  );
  assign axi_ar_ready = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_r_valid = 3'h2 == state; // @[Mux.scala 81:61]
  assign axi_r_bits_data = RamBB_i1_rdata; // @[sram_AxiLite.scala 98:21]
  assign axi_aw_ready = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_w_ready = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_b_valid = 3'h4 == state; // @[Mux.scala 81:61]
  assign RamBB_i1_clock = clock; // @[sram_AxiLite.scala 78:25]
  assign RamBB_i1_addr = _T_8 ? axi_aw_bits_addr : _RamBB_i1_io_addr_T_1; // @[Mux.scala 81:58]
  assign RamBB_i1_mem_wen = 3'h4 == state; // @[Mux.scala 81:61]
  assign RamBB_i1_valid = _T_8 | _T_6; // @[Mux.scala 81:58]
  assign RamBB_i1_wdata = axi_w_bits_data; // @[sram_AxiLite.scala 92:25]
  assign RamBB_i1_wmask = axi_w_bits_strb; // @[sram_AxiLite.scala 93:25]
  always @(posedge clock) begin
    if (reset) begin // @[sram_AxiLite.scala 42:24]
      delay <= 1'h0; // @[sram_AxiLite.scala 42:24]
    end else if (3'h0 == state) begin // @[sram_AxiLite.scala 47:20]
      delay <= 1'h0; // @[sram_AxiLite.scala 49:19]
    end else if (3'h1 == state) begin // @[sram_AxiLite.scala 47:20]
      delay <= delay - 1'h1; // @[sram_AxiLite.scala 63:19]
    end else if (!(3'h2 == state)) begin // @[sram_AxiLite.scala 47:20]
      delay <= _GEN_4;
    end
    if (reset) begin // @[sram_AxiLite.scala 46:24]
      state <= 3'h0; // @[sram_AxiLite.scala 46:24]
    end else if (3'h0 == state) begin // @[sram_AxiLite.scala 47:20]
      if (_T_1) begin // @[sram_AxiLite.scala 51:32]
        state <= 3'h1; // @[sram_AxiLite.scala 52:23]
      end else if (_T_2 & _T_3) begin // @[sram_AxiLite.scala 54:51]
        state <= 3'h3; // @[sram_AxiLite.scala 55:23]
      end else begin
        state <= 3'h0; // @[sram_AxiLite.scala 58:23]
      end
    end else if (3'h1 == state) begin // @[sram_AxiLite.scala 47:20]
      if (~delay) begin // @[sram_AxiLite.scala 62:25]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[sram_AxiLite.scala 47:20]
      state <= _state_T_3; // @[sram_AxiLite.scala 66:19]
    end else begin
      state <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_out_inst,
  output [31:0] io_out_pc,
  output [31:0] io_out_difftest_mcause,
  output [31:0] io_out_difftest_mepc,
  output [31:0] io_out_difftest_mstatus,
  output [31:0] io_out_difftest_mtvec,
  output        io_out_wb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  IDU_i_from_IFU_valid; // @[core.scala 32:27]
  wire [31:0] IDU_i_from_IFU_bits_inst; // @[core.scala 32:27]
  wire [31:0] IDU_i_from_IFU_bits_pc; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_valid; // @[core.scala 32:27]
  wire [31:0] IDU_i_to_ISU_bits_imm; // @[core.scala 32:27]
  wire [31:0] IDU_i_to_ISU_bits_pc; // @[core.scala 32:27]
  wire [4:0] IDU_i_to_ISU_bits_rs1; // @[core.scala 32:27]
  wire [4:0] IDU_i_to_ISU_bits_rs2; // @[core.scala 32:27]
  wire [4:0] IDU_i_to_ISU_bits_rd; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_reg_wen; // @[core.scala 32:27]
  wire [2:0] IDU_i_to_ISU_bits_ctrl_sig_fu_op; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_mem_wen; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_is_ebreak; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_not_impl; // @[core.scala 32:27]
  wire [1:0] IDU_i_to_ISU_bits_ctrl_sig_src1_op; // @[core.scala 32:27]
  wire [1:0] IDU_i_to_ISU_bits_ctrl_sig_src2_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_alu_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_lsu_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_bru_op; // @[core.scala 32:27]
  wire [2:0] IDU_i_to_ISU_bits_ctrl_sig_csr_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_mdu_op; // @[core.scala 32:27]
  wire  ISU_i_clock; // @[core.scala 33:27]
  wire  ISU_i_reset; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_valid; // @[core.scala 33:27]
  wire [31:0] ISU_i_from_IDU_bits_imm; // @[core.scala 33:27]
  wire [31:0] ISU_i_from_IDU_bits_pc; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_IDU_bits_rs1; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_IDU_bits_rs2; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_IDU_bits_rd; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_reg_wen; // @[core.scala 33:27]
  wire [2:0] ISU_i_from_IDU_bits_ctrl_sig_fu_op; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_mem_wen; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_is_ebreak; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_not_impl; // @[core.scala 33:27]
  wire [1:0] ISU_i_from_IDU_bits_ctrl_sig_src1_op; // @[core.scala 33:27]
  wire [1:0] ISU_i_from_IDU_bits_ctrl_sig_src2_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_alu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_lsu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_bru_op; // @[core.scala 33:27]
  wire [2:0] ISU_i_from_IDU_bits_ctrl_sig_csr_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_mdu_op; // @[core.scala 33:27]
  wire  ISU_i_from_WBU_bits_reg_wen; // @[core.scala 33:27]
  wire [31:0] ISU_i_from_WBU_bits_wdata; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_WBU_bits_rd; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_valid; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_imm; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_pc; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_rdata1; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_rdata2; // @[core.scala 33:27]
  wire [4:0] ISU_i_to_EXU_bits_rd; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_reg_wen; // @[core.scala 33:27]
  wire [2:0] ISU_i_to_EXU_bits_ctrl_sig_fu_op; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_mem_wen; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_is_ebreak; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_not_impl; // @[core.scala 33:27]
  wire [1:0] ISU_i_to_EXU_bits_ctrl_sig_src1_op; // @[core.scala 33:27]
  wire [1:0] ISU_i_to_EXU_bits_ctrl_sig_src2_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_alu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_lsu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_bru_op; // @[core.scala 33:27]
  wire [2:0] ISU_i_to_EXU_bits_ctrl_sig_csr_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_mdu_op; // @[core.scala 33:27]
  wire  EXU_i_clock; // @[core.scala 34:27]
  wire  EXU_i_reset; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_ready; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_imm; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_pc; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_rdata1; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_rdata2; // @[core.scala 34:27]
  wire [4:0] EXU_i_from_ISU_bits_rd; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_reg_wen; // @[core.scala 34:27]
  wire [2:0] EXU_i_from_ISU_bits_ctrl_sig_fu_op; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_mem_wen; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_is_ebreak; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_not_impl; // @[core.scala 34:27]
  wire [1:0] EXU_i_from_ISU_bits_ctrl_sig_src1_op; // @[core.scala 34:27]
  wire [1:0] EXU_i_from_ISU_bits_ctrl_sig_src2_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_alu_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_lsu_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_bru_op; // @[core.scala 34:27]
  wire [2:0] EXU_i_from_ISU_bits_ctrl_sig_csr_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_mdu_op; // @[core.scala 34:27]
  wire  EXU_i_to_WBU_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_alu_result; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_mdu_result; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_lsu_rdata; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_csr_rdata; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_pc; // @[core.scala 34:27]
  wire  EXU_i_to_WBU_bits_reg_wen; // @[core.scala 34:27]
  wire [4:0] EXU_i_to_WBU_bits_rd; // @[core.scala 34:27]
  wire [2:0] EXU_i_to_WBU_bits_fu_op; // @[core.scala 34:27]
  wire  EXU_i_to_IFU_bits_bru_ctrl_br; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_IFU_bits_bru_addr; // @[core.scala 34:27]
  wire  EXU_i_to_IFU_bits_csr_ctrl_br; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_IFU_bits_csr_addr; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mcause; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mepc; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mstatus; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mtvec; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_ar_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_ar_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_ar_bits_addr; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_r_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_r_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_r_bits_data; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_aw_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_aw_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_aw_bits_addr; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_w_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_w_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_w_bits_data; // @[core.scala 34:27]
  wire [3:0] EXU_i_lsu_axi_master_w_bits_strb; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_b_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_b_valid; // @[core.scala 34:27]
  wire  WBU_i_from_EXU_ready; // @[core.scala 35:27]
  wire  WBU_i_from_EXU_valid; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_alu_result; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_mdu_result; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_lsu_rdata; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_csr_rdata; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_pc; // @[core.scala 35:27]
  wire  WBU_i_from_EXU_bits_reg_wen; // @[core.scala 35:27]
  wire [4:0] WBU_i_from_EXU_bits_rd; // @[core.scala 35:27]
  wire [2:0] WBU_i_from_EXU_bits_fu_op; // @[core.scala 35:27]
  wire  WBU_i_to_ISU_bits_reg_wen; // @[core.scala 35:27]
  wire [31:0] WBU_i_to_ISU_bits_wdata; // @[core.scala 35:27]
  wire [4:0] WBU_i_to_ISU_bits_rd; // @[core.scala 35:27]
  wire  WBU_i_to_IFU_valid; // @[core.scala 35:27]
  wire  IFU_i_clock; // @[core.scala 48:27]
  wire  IFU_i_reset; // @[core.scala 48:27]
  wire  IFU_i_to_IDU_valid; // @[core.scala 48:27]
  wire [31:0] IFU_i_to_IDU_bits_inst; // @[core.scala 48:27]
  wire [31:0] IFU_i_to_IDU_bits_pc; // @[core.scala 48:27]
  wire  IFU_i_from_EXU_bits_bru_ctrl_br; // @[core.scala 48:27]
  wire [31:0] IFU_i_from_EXU_bits_bru_addr; // @[core.scala 48:27]
  wire  IFU_i_from_EXU_bits_csr_ctrl_br; // @[core.scala 48:27]
  wire [31:0] IFU_i_from_EXU_bits_csr_addr; // @[core.scala 48:27]
  wire  IFU_i_from_WBU_ready; // @[core.scala 48:27]
  wire  IFU_i_from_WBU_valid; // @[core.scala 48:27]
  wire  IFU_i_to_cache_ready; // @[core.scala 48:27]
  wire  IFU_i_to_cache_valid; // @[core.scala 48:27]
  wire [31:0] IFU_i_to_cache_bits_addr; // @[core.scala 48:27]
  wire  IFU_i_from_cache_ready; // @[core.scala 48:27]
  wire  IFU_i_from_cache_valid; // @[core.scala 48:27]
  wire [31:0] IFU_i_from_cache_bits_data; // @[core.scala 48:27]
  wire  icache_clock; // @[core.scala 49:27]
  wire  icache_reset; // @[core.scala 49:27]
  wire  icache_from_IFU_ready; // @[core.scala 49:27]
  wire  icache_from_IFU_valid; // @[core.scala 49:27]
  wire [31:0] icache_from_IFU_bits_addr; // @[core.scala 49:27]
  wire  icache_to_IFU_valid; // @[core.scala 49:27]
  wire [31:0] icache_to_IFU_bits_data; // @[core.scala 49:27]
  wire  icache_to_sram_ar_ready; // @[core.scala 49:27]
  wire  icache_to_sram_ar_valid; // @[core.scala 49:27]
  wire [31:0] icache_to_sram_ar_bits_addr; // @[core.scala 49:27]
  wire [7:0] icache_to_sram_ar_bits_len; // @[core.scala 49:27]
  wire  icache_to_sram_r_ready; // @[core.scala 49:27]
  wire  icache_to_sram_r_valid; // @[core.scala 49:27]
  wire [31:0] icache_to_sram_r_bits_data; // @[core.scala 49:27]
  wire  icache_to_sram_r_bits_last; // @[core.scala 49:27]
  wire  sram_i_clock; // @[core.scala 50:27]
  wire  sram_i_reset; // @[core.scala 50:27]
  wire  sram_i_axi_ar_ready; // @[core.scala 50:27]
  wire  sram_i_axi_ar_valid; // @[core.scala 50:27]
  wire [31:0] sram_i_axi_ar_bits_addr; // @[core.scala 50:27]
  wire [7:0] sram_i_axi_ar_bits_len; // @[core.scala 50:27]
  wire  sram_i_axi_r_ready; // @[core.scala 50:27]
  wire  sram_i_axi_r_valid; // @[core.scala 50:27]
  wire [31:0] sram_i_axi_r_bits_data; // @[core.scala 50:27]
  wire  sram_i_axi_r_bits_last; // @[core.scala 50:27]
  wire  sram_i2_clock; // @[core.scala 57:27]
  wire  sram_i2_reset; // @[core.scala 57:27]
  wire  sram_i2_axi_ar_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_ar_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_ar_bits_addr; // @[core.scala 57:27]
  wire  sram_i2_axi_r_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_r_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_r_bits_data; // @[core.scala 57:27]
  wire  sram_i2_axi_aw_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_aw_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_aw_bits_addr; // @[core.scala 57:27]
  wire  sram_i2_axi_w_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_w_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_w_bits_data; // @[core.scala 57:27]
  wire [3:0] sram_i2_axi_w_bits_strb; // @[core.scala 57:27]
  wire  sram_i2_axi_b_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_b_valid; // @[core.scala 57:27]
  wire  _EXU_i_from_ISU_bits_T = ISU_i_to_EXU_valid & EXU_i_from_ISU_ready; // @[Connect.scala 26:58]
  reg [31:0] EXU_i_from_ISU_bits_r_imm; // @[Reg.scala 19:16]
  reg [31:0] EXU_i_from_ISU_bits_r_pc; // @[Reg.scala 19:16]
  reg [31:0] EXU_i_from_ISU_bits_r_rdata1; // @[Reg.scala 19:16]
  reg [31:0] EXU_i_from_ISU_bits_r_rdata2; // @[Reg.scala 19:16]
  reg [4:0] EXU_i_from_ISU_bits_r_rd; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen; // @[Reg.scala 19:16]
  reg [2:0] EXU_i_from_ISU_bits_r_ctrl_sig_fu_op; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_not_impl; // @[Reg.scala 19:16]
  reg [1:0] EXU_i_from_ISU_bits_r_ctrl_sig_src1_op; // @[Reg.scala 19:16]
  reg [1:0] EXU_i_from_ISU_bits_r_ctrl_sig_src2_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_alu_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_bru_op; // @[Reg.scala 19:16]
  reg [2:0] EXU_i_from_ISU_bits_r_ctrl_sig_csr_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op; // @[Reg.scala 19:16]
  IDU IDU_i ( // @[core.scala 32:27]
    .from_IFU_valid(IDU_i_from_IFU_valid),
    .from_IFU_bits_inst(IDU_i_from_IFU_bits_inst),
    .from_IFU_bits_pc(IDU_i_from_IFU_bits_pc),
    .to_ISU_valid(IDU_i_to_ISU_valid),
    .to_ISU_bits_imm(IDU_i_to_ISU_bits_imm),
    .to_ISU_bits_pc(IDU_i_to_ISU_bits_pc),
    .to_ISU_bits_rs1(IDU_i_to_ISU_bits_rs1),
    .to_ISU_bits_rs2(IDU_i_to_ISU_bits_rs2),
    .to_ISU_bits_rd(IDU_i_to_ISU_bits_rd),
    .to_ISU_bits_ctrl_sig_reg_wen(IDU_i_to_ISU_bits_ctrl_sig_reg_wen),
    .to_ISU_bits_ctrl_sig_fu_op(IDU_i_to_ISU_bits_ctrl_sig_fu_op),
    .to_ISU_bits_ctrl_sig_mem_wen(IDU_i_to_ISU_bits_ctrl_sig_mem_wen),
    .to_ISU_bits_ctrl_sig_is_ebreak(IDU_i_to_ISU_bits_ctrl_sig_is_ebreak),
    .to_ISU_bits_ctrl_sig_not_impl(IDU_i_to_ISU_bits_ctrl_sig_not_impl),
    .to_ISU_bits_ctrl_sig_src1_op(IDU_i_to_ISU_bits_ctrl_sig_src1_op),
    .to_ISU_bits_ctrl_sig_src2_op(IDU_i_to_ISU_bits_ctrl_sig_src2_op),
    .to_ISU_bits_ctrl_sig_alu_op(IDU_i_to_ISU_bits_ctrl_sig_alu_op),
    .to_ISU_bits_ctrl_sig_lsu_op(IDU_i_to_ISU_bits_ctrl_sig_lsu_op),
    .to_ISU_bits_ctrl_sig_bru_op(IDU_i_to_ISU_bits_ctrl_sig_bru_op),
    .to_ISU_bits_ctrl_sig_csr_op(IDU_i_to_ISU_bits_ctrl_sig_csr_op),
    .to_ISU_bits_ctrl_sig_mdu_op(IDU_i_to_ISU_bits_ctrl_sig_mdu_op)
  );
  ISU ISU_i ( // @[core.scala 33:27]
    .clock(ISU_i_clock),
    .reset(ISU_i_reset),
    .from_IDU_valid(ISU_i_from_IDU_valid),
    .from_IDU_bits_imm(ISU_i_from_IDU_bits_imm),
    .from_IDU_bits_pc(ISU_i_from_IDU_bits_pc),
    .from_IDU_bits_rs1(ISU_i_from_IDU_bits_rs1),
    .from_IDU_bits_rs2(ISU_i_from_IDU_bits_rs2),
    .from_IDU_bits_rd(ISU_i_from_IDU_bits_rd),
    .from_IDU_bits_ctrl_sig_reg_wen(ISU_i_from_IDU_bits_ctrl_sig_reg_wen),
    .from_IDU_bits_ctrl_sig_fu_op(ISU_i_from_IDU_bits_ctrl_sig_fu_op),
    .from_IDU_bits_ctrl_sig_mem_wen(ISU_i_from_IDU_bits_ctrl_sig_mem_wen),
    .from_IDU_bits_ctrl_sig_is_ebreak(ISU_i_from_IDU_bits_ctrl_sig_is_ebreak),
    .from_IDU_bits_ctrl_sig_not_impl(ISU_i_from_IDU_bits_ctrl_sig_not_impl),
    .from_IDU_bits_ctrl_sig_src1_op(ISU_i_from_IDU_bits_ctrl_sig_src1_op),
    .from_IDU_bits_ctrl_sig_src2_op(ISU_i_from_IDU_bits_ctrl_sig_src2_op),
    .from_IDU_bits_ctrl_sig_alu_op(ISU_i_from_IDU_bits_ctrl_sig_alu_op),
    .from_IDU_bits_ctrl_sig_lsu_op(ISU_i_from_IDU_bits_ctrl_sig_lsu_op),
    .from_IDU_bits_ctrl_sig_bru_op(ISU_i_from_IDU_bits_ctrl_sig_bru_op),
    .from_IDU_bits_ctrl_sig_csr_op(ISU_i_from_IDU_bits_ctrl_sig_csr_op),
    .from_IDU_bits_ctrl_sig_mdu_op(ISU_i_from_IDU_bits_ctrl_sig_mdu_op),
    .from_WBU_bits_reg_wen(ISU_i_from_WBU_bits_reg_wen),
    .from_WBU_bits_wdata(ISU_i_from_WBU_bits_wdata),
    .from_WBU_bits_rd(ISU_i_from_WBU_bits_rd),
    .to_EXU_valid(ISU_i_to_EXU_valid),
    .to_EXU_bits_imm(ISU_i_to_EXU_bits_imm),
    .to_EXU_bits_pc(ISU_i_to_EXU_bits_pc),
    .to_EXU_bits_rdata1(ISU_i_to_EXU_bits_rdata1),
    .to_EXU_bits_rdata2(ISU_i_to_EXU_bits_rdata2),
    .to_EXU_bits_rd(ISU_i_to_EXU_bits_rd),
    .to_EXU_bits_ctrl_sig_reg_wen(ISU_i_to_EXU_bits_ctrl_sig_reg_wen),
    .to_EXU_bits_ctrl_sig_fu_op(ISU_i_to_EXU_bits_ctrl_sig_fu_op),
    .to_EXU_bits_ctrl_sig_mem_wen(ISU_i_to_EXU_bits_ctrl_sig_mem_wen),
    .to_EXU_bits_ctrl_sig_is_ebreak(ISU_i_to_EXU_bits_ctrl_sig_is_ebreak),
    .to_EXU_bits_ctrl_sig_not_impl(ISU_i_to_EXU_bits_ctrl_sig_not_impl),
    .to_EXU_bits_ctrl_sig_src1_op(ISU_i_to_EXU_bits_ctrl_sig_src1_op),
    .to_EXU_bits_ctrl_sig_src2_op(ISU_i_to_EXU_bits_ctrl_sig_src2_op),
    .to_EXU_bits_ctrl_sig_alu_op(ISU_i_to_EXU_bits_ctrl_sig_alu_op),
    .to_EXU_bits_ctrl_sig_lsu_op(ISU_i_to_EXU_bits_ctrl_sig_lsu_op),
    .to_EXU_bits_ctrl_sig_bru_op(ISU_i_to_EXU_bits_ctrl_sig_bru_op),
    .to_EXU_bits_ctrl_sig_csr_op(ISU_i_to_EXU_bits_ctrl_sig_csr_op),
    .to_EXU_bits_ctrl_sig_mdu_op(ISU_i_to_EXU_bits_ctrl_sig_mdu_op)
  );
  EXU EXU_i ( // @[core.scala 34:27]
    .clock(EXU_i_clock),
    .reset(EXU_i_reset),
    .from_ISU_ready(EXU_i_from_ISU_ready),
    .from_ISU_valid(EXU_i_from_ISU_valid),
    .from_ISU_bits_imm(EXU_i_from_ISU_bits_imm),
    .from_ISU_bits_pc(EXU_i_from_ISU_bits_pc),
    .from_ISU_bits_rdata1(EXU_i_from_ISU_bits_rdata1),
    .from_ISU_bits_rdata2(EXU_i_from_ISU_bits_rdata2),
    .from_ISU_bits_rd(EXU_i_from_ISU_bits_rd),
    .from_ISU_bits_ctrl_sig_reg_wen(EXU_i_from_ISU_bits_ctrl_sig_reg_wen),
    .from_ISU_bits_ctrl_sig_fu_op(EXU_i_from_ISU_bits_ctrl_sig_fu_op),
    .from_ISU_bits_ctrl_sig_mem_wen(EXU_i_from_ISU_bits_ctrl_sig_mem_wen),
    .from_ISU_bits_ctrl_sig_is_ebreak(EXU_i_from_ISU_bits_ctrl_sig_is_ebreak),
    .from_ISU_bits_ctrl_sig_not_impl(EXU_i_from_ISU_bits_ctrl_sig_not_impl),
    .from_ISU_bits_ctrl_sig_src1_op(EXU_i_from_ISU_bits_ctrl_sig_src1_op),
    .from_ISU_bits_ctrl_sig_src2_op(EXU_i_from_ISU_bits_ctrl_sig_src2_op),
    .from_ISU_bits_ctrl_sig_alu_op(EXU_i_from_ISU_bits_ctrl_sig_alu_op),
    .from_ISU_bits_ctrl_sig_lsu_op(EXU_i_from_ISU_bits_ctrl_sig_lsu_op),
    .from_ISU_bits_ctrl_sig_bru_op(EXU_i_from_ISU_bits_ctrl_sig_bru_op),
    .from_ISU_bits_ctrl_sig_csr_op(EXU_i_from_ISU_bits_ctrl_sig_csr_op),
    .from_ISU_bits_ctrl_sig_mdu_op(EXU_i_from_ISU_bits_ctrl_sig_mdu_op),
    .to_WBU_valid(EXU_i_to_WBU_valid),
    .to_WBU_bits_alu_result(EXU_i_to_WBU_bits_alu_result),
    .to_WBU_bits_mdu_result(EXU_i_to_WBU_bits_mdu_result),
    .to_WBU_bits_lsu_rdata(EXU_i_to_WBU_bits_lsu_rdata),
    .to_WBU_bits_csr_rdata(EXU_i_to_WBU_bits_csr_rdata),
    .to_WBU_bits_pc(EXU_i_to_WBU_bits_pc),
    .to_WBU_bits_reg_wen(EXU_i_to_WBU_bits_reg_wen),
    .to_WBU_bits_rd(EXU_i_to_WBU_bits_rd),
    .to_WBU_bits_fu_op(EXU_i_to_WBU_bits_fu_op),
    .to_IFU_bits_bru_ctrl_br(EXU_i_to_IFU_bits_bru_ctrl_br),
    .to_IFU_bits_bru_addr(EXU_i_to_IFU_bits_bru_addr),
    .to_IFU_bits_csr_ctrl_br(EXU_i_to_IFU_bits_csr_ctrl_br),
    .to_IFU_bits_csr_addr(EXU_i_to_IFU_bits_csr_addr),
    .difftest_mcause(EXU_i_difftest_mcause),
    .difftest_mepc(EXU_i_difftest_mepc),
    .difftest_mstatus(EXU_i_difftest_mstatus),
    .difftest_mtvec(EXU_i_difftest_mtvec),
    .lsu_axi_master_ar_ready(EXU_i_lsu_axi_master_ar_ready),
    .lsu_axi_master_ar_valid(EXU_i_lsu_axi_master_ar_valid),
    .lsu_axi_master_ar_bits_addr(EXU_i_lsu_axi_master_ar_bits_addr),
    .lsu_axi_master_r_ready(EXU_i_lsu_axi_master_r_ready),
    .lsu_axi_master_r_valid(EXU_i_lsu_axi_master_r_valid),
    .lsu_axi_master_r_bits_data(EXU_i_lsu_axi_master_r_bits_data),
    .lsu_axi_master_aw_ready(EXU_i_lsu_axi_master_aw_ready),
    .lsu_axi_master_aw_valid(EXU_i_lsu_axi_master_aw_valid),
    .lsu_axi_master_aw_bits_addr(EXU_i_lsu_axi_master_aw_bits_addr),
    .lsu_axi_master_w_ready(EXU_i_lsu_axi_master_w_ready),
    .lsu_axi_master_w_valid(EXU_i_lsu_axi_master_w_valid),
    .lsu_axi_master_w_bits_data(EXU_i_lsu_axi_master_w_bits_data),
    .lsu_axi_master_w_bits_strb(EXU_i_lsu_axi_master_w_bits_strb),
    .lsu_axi_master_b_ready(EXU_i_lsu_axi_master_b_ready),
    .lsu_axi_master_b_valid(EXU_i_lsu_axi_master_b_valid)
  );
  WBU WBU_i ( // @[core.scala 35:27]
    .from_EXU_ready(WBU_i_from_EXU_ready),
    .from_EXU_valid(WBU_i_from_EXU_valid),
    .from_EXU_bits_alu_result(WBU_i_from_EXU_bits_alu_result),
    .from_EXU_bits_mdu_result(WBU_i_from_EXU_bits_mdu_result),
    .from_EXU_bits_lsu_rdata(WBU_i_from_EXU_bits_lsu_rdata),
    .from_EXU_bits_csr_rdata(WBU_i_from_EXU_bits_csr_rdata),
    .from_EXU_bits_pc(WBU_i_from_EXU_bits_pc),
    .from_EXU_bits_reg_wen(WBU_i_from_EXU_bits_reg_wen),
    .from_EXU_bits_rd(WBU_i_from_EXU_bits_rd),
    .from_EXU_bits_fu_op(WBU_i_from_EXU_bits_fu_op),
    .to_ISU_bits_reg_wen(WBU_i_to_ISU_bits_reg_wen),
    .to_ISU_bits_wdata(WBU_i_to_ISU_bits_wdata),
    .to_ISU_bits_rd(WBU_i_to_ISU_bits_rd),
    .to_IFU_valid(WBU_i_to_IFU_valid)
  );
  IFU_cache IFU_i ( // @[core.scala 48:27]
    .clock(IFU_i_clock),
    .reset(IFU_i_reset),
    .to_IDU_valid(IFU_i_to_IDU_valid),
    .to_IDU_bits_inst(IFU_i_to_IDU_bits_inst),
    .to_IDU_bits_pc(IFU_i_to_IDU_bits_pc),
    .from_EXU_bits_bru_ctrl_br(IFU_i_from_EXU_bits_bru_ctrl_br),
    .from_EXU_bits_bru_addr(IFU_i_from_EXU_bits_bru_addr),
    .from_EXU_bits_csr_ctrl_br(IFU_i_from_EXU_bits_csr_ctrl_br),
    .from_EXU_bits_csr_addr(IFU_i_from_EXU_bits_csr_addr),
    .from_WBU_ready(IFU_i_from_WBU_ready),
    .from_WBU_valid(IFU_i_from_WBU_valid),
    .to_cache_ready(IFU_i_to_cache_ready),
    .to_cache_valid(IFU_i_to_cache_valid),
    .to_cache_bits_addr(IFU_i_to_cache_bits_addr),
    .from_cache_ready(IFU_i_from_cache_ready),
    .from_cache_valid(IFU_i_from_cache_valid),
    .from_cache_bits_data(IFU_i_from_cache_bits_data)
  );
  I_Cache icache ( // @[core.scala 49:27]
    .clock(icache_clock),
    .reset(icache_reset),
    .from_IFU_ready(icache_from_IFU_ready),
    .from_IFU_valid(icache_from_IFU_valid),
    .from_IFU_bits_addr(icache_from_IFU_bits_addr),
    .to_IFU_valid(icache_to_IFU_valid),
    .to_IFU_bits_data(icache_to_IFU_bits_data),
    .to_sram_ar_ready(icache_to_sram_ar_ready),
    .to_sram_ar_valid(icache_to_sram_ar_valid),
    .to_sram_ar_bits_addr(icache_to_sram_ar_bits_addr),
    .to_sram_ar_bits_len(icache_to_sram_ar_bits_len),
    .to_sram_r_ready(icache_to_sram_r_ready),
    .to_sram_r_valid(icache_to_sram_r_valid),
    .to_sram_r_bits_data(icache_to_sram_r_bits_data),
    .to_sram_r_bits_last(icache_to_sram_r_bits_last)
  );
  SRAM_axi sram_i ( // @[core.scala 50:27]
    .clock(sram_i_clock),
    .reset(sram_i_reset),
    .axi_ar_ready(sram_i_axi_ar_ready),
    .axi_ar_valid(sram_i_axi_ar_valid),
    .axi_ar_bits_addr(sram_i_axi_ar_bits_addr),
    .axi_ar_bits_len(sram_i_axi_ar_bits_len),
    .axi_r_ready(sram_i_axi_r_ready),
    .axi_r_valid(sram_i_axi_r_valid),
    .axi_r_bits_data(sram_i_axi_r_bits_data),
    .axi_r_bits_last(sram_i_axi_r_bits_last)
  );
  SRAM sram_i2 ( // @[core.scala 57:27]
    .clock(sram_i2_clock),
    .reset(sram_i2_reset),
    .axi_ar_ready(sram_i2_axi_ar_ready),
    .axi_ar_valid(sram_i2_axi_ar_valid),
    .axi_ar_bits_addr(sram_i2_axi_ar_bits_addr),
    .axi_r_ready(sram_i2_axi_r_ready),
    .axi_r_valid(sram_i2_axi_r_valid),
    .axi_r_bits_data(sram_i2_axi_r_bits_data),
    .axi_aw_ready(sram_i2_axi_aw_ready),
    .axi_aw_valid(sram_i2_axi_aw_valid),
    .axi_aw_bits_addr(sram_i2_axi_aw_bits_addr),
    .axi_w_ready(sram_i2_axi_w_ready),
    .axi_w_valid(sram_i2_axi_w_valid),
    .axi_w_bits_data(sram_i2_axi_w_bits_data),
    .axi_w_bits_strb(sram_i2_axi_w_bits_strb),
    .axi_b_ready(sram_i2_axi_b_ready),
    .axi_b_valid(sram_i2_axi_b_valid)
  );
  assign io_out_inst = IFU_i_to_IDU_bits_inst; // @[core.scala 75:20]
  assign io_out_pc = IFU_i_to_IDU_bits_pc; // @[core.scala 76:20]
  assign io_out_difftest_mcause = EXU_i_difftest_mcause; // @[core.scala 79:21]
  assign io_out_difftest_mepc = EXU_i_difftest_mepc; // @[core.scala 79:21]
  assign io_out_difftest_mstatus = EXU_i_difftest_mstatus; // @[core.scala 79:21]
  assign io_out_difftest_mtvec = EXU_i_difftest_mtvec; // @[core.scala 79:21]
  assign io_out_wb = WBU_i_to_IFU_valid; // @[core.scala 77:20]
  assign IDU_i_from_IFU_valid = IFU_i_to_IDU_valid; // @[Connect.scala 16:22]
  assign IDU_i_from_IFU_bits_inst = IFU_i_to_IDU_bits_inst; // @[Connect.scala 15:22]
  assign IDU_i_from_IFU_bits_pc = IFU_i_to_IDU_bits_pc; // @[Connect.scala 15:22]
  assign ISU_i_clock = clock;
  assign ISU_i_reset = reset;
  assign ISU_i_from_IDU_valid = IDU_i_to_ISU_valid; // @[Connect.scala 16:22]
  assign ISU_i_from_IDU_bits_imm = IDU_i_to_ISU_bits_imm; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_pc = IDU_i_to_ISU_bits_pc; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_rs1 = IDU_i_to_ISU_bits_rs1; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_rs2 = IDU_i_to_ISU_bits_rs2; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_rd = IDU_i_to_ISU_bits_rd; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_reg_wen = IDU_i_to_ISU_bits_ctrl_sig_reg_wen; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_fu_op = IDU_i_to_ISU_bits_ctrl_sig_fu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_mem_wen = IDU_i_to_ISU_bits_ctrl_sig_mem_wen; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_is_ebreak = IDU_i_to_ISU_bits_ctrl_sig_is_ebreak; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_not_impl = IDU_i_to_ISU_bits_ctrl_sig_not_impl; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_src1_op = IDU_i_to_ISU_bits_ctrl_sig_src1_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_src2_op = IDU_i_to_ISU_bits_ctrl_sig_src2_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_alu_op = IDU_i_to_ISU_bits_ctrl_sig_alu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_lsu_op = IDU_i_to_ISU_bits_ctrl_sig_lsu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_bru_op = IDU_i_to_ISU_bits_ctrl_sig_bru_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_csr_op = IDU_i_to_ISU_bits_ctrl_sig_csr_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_mdu_op = IDU_i_to_ISU_bits_ctrl_sig_mdu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_WBU_bits_reg_wen = WBU_i_to_ISU_bits_reg_wen; // @[Connect.scala 15:22]
  assign ISU_i_from_WBU_bits_wdata = WBU_i_to_ISU_bits_wdata; // @[Connect.scala 15:22]
  assign ISU_i_from_WBU_bits_rd = WBU_i_to_ISU_bits_rd; // @[Connect.scala 15:22]
  assign EXU_i_clock = clock;
  assign EXU_i_reset = reset;
  assign EXU_i_from_ISU_valid = ISU_i_to_EXU_valid; // @[Connect.scala 27:22]
  assign EXU_i_from_ISU_bits_imm = EXU_i_from_ISU_bits_r_imm; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_pc = EXU_i_from_ISU_bits_r_pc; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_rdata1 = EXU_i_from_ISU_bits_r_rdata1; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_rdata2 = EXU_i_from_ISU_bits_r_rdata2; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_rd = EXU_i_from_ISU_bits_r_rd; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_reg_wen = EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_fu_op = EXU_i_from_ISU_bits_r_ctrl_sig_fu_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_mem_wen = EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_is_ebreak = EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_not_impl = EXU_i_from_ISU_bits_r_ctrl_sig_not_impl; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_src1_op = EXU_i_from_ISU_bits_r_ctrl_sig_src1_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_src2_op = EXU_i_from_ISU_bits_r_ctrl_sig_src2_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_alu_op = EXU_i_from_ISU_bits_r_ctrl_sig_alu_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_lsu_op = EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_bru_op = EXU_i_from_ISU_bits_r_ctrl_sig_bru_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_csr_op = EXU_i_from_ISU_bits_r_ctrl_sig_csr_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_mdu_op = EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op; // @[Connect.scala 26:22]
  assign EXU_i_lsu_axi_master_ar_ready = sram_i2_axi_ar_ready; // @[Connect.scala 17:22]
  assign EXU_i_lsu_axi_master_r_valid = sram_i2_axi_r_valid; // @[Connect.scala 16:22]
  assign EXU_i_lsu_axi_master_r_bits_data = sram_i2_axi_r_bits_data; // @[Connect.scala 15:22]
  assign EXU_i_lsu_axi_master_aw_ready = sram_i2_axi_aw_ready; // @[Connect.scala 17:22]
  assign EXU_i_lsu_axi_master_w_ready = sram_i2_axi_w_ready; // @[Connect.scala 17:22]
  assign EXU_i_lsu_axi_master_b_valid = sram_i2_axi_b_valid; // @[Connect.scala 16:22]
  assign WBU_i_from_EXU_valid = EXU_i_to_WBU_valid; // @[Connect.scala 16:22]
  assign WBU_i_from_EXU_bits_alu_result = EXU_i_to_WBU_bits_alu_result; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_mdu_result = EXU_i_to_WBU_bits_mdu_result; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_lsu_rdata = EXU_i_to_WBU_bits_lsu_rdata; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_csr_rdata = EXU_i_to_WBU_bits_csr_rdata; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_pc = EXU_i_to_WBU_bits_pc; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_reg_wen = EXU_i_to_WBU_bits_reg_wen; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_rd = EXU_i_to_WBU_bits_rd; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_fu_op = EXU_i_to_WBU_bits_fu_op; // @[Connect.scala 15:22]
  assign IFU_i_clock = clock;
  assign IFU_i_reset = reset;
  assign IFU_i_from_EXU_bits_bru_ctrl_br = EXU_i_to_IFU_bits_bru_ctrl_br; // @[Connect.scala 15:22]
  assign IFU_i_from_EXU_bits_bru_addr = EXU_i_to_IFU_bits_bru_addr; // @[Connect.scala 15:22]
  assign IFU_i_from_EXU_bits_csr_ctrl_br = EXU_i_to_IFU_bits_csr_ctrl_br; // @[Connect.scala 15:22]
  assign IFU_i_from_EXU_bits_csr_addr = EXU_i_to_IFU_bits_csr_addr; // @[Connect.scala 15:22]
  assign IFU_i_from_WBU_valid = WBU_i_to_IFU_valid; // @[Connect.scala 16:22]
  assign IFU_i_to_cache_ready = icache_from_IFU_ready; // @[Connect.scala 17:22]
  assign IFU_i_from_cache_valid = icache_to_IFU_valid; // @[Connect.scala 16:22]
  assign IFU_i_from_cache_bits_data = icache_to_IFU_bits_data; // @[Connect.scala 15:22]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_from_IFU_valid = IFU_i_to_cache_valid; // @[Connect.scala 16:22]
  assign icache_from_IFU_bits_addr = IFU_i_to_cache_bits_addr; // @[Connect.scala 15:22]
  assign icache_to_sram_ar_ready = sram_i_axi_ar_ready; // @[Connect.scala 17:22]
  assign icache_to_sram_r_valid = sram_i_axi_r_valid; // @[Connect.scala 16:22]
  assign icache_to_sram_r_bits_data = sram_i_axi_r_bits_data; // @[Connect.scala 15:22]
  assign icache_to_sram_r_bits_last = sram_i_axi_r_bits_last; // @[Connect.scala 15:22]
  assign sram_i_clock = clock;
  assign sram_i_reset = reset;
  assign sram_i_axi_ar_valid = icache_to_sram_ar_valid; // @[Connect.scala 16:22]
  assign sram_i_axi_ar_bits_addr = icache_to_sram_ar_bits_addr; // @[Connect.scala 15:22]
  assign sram_i_axi_ar_bits_len = icache_to_sram_ar_bits_len; // @[Connect.scala 15:22]
  assign sram_i_axi_r_ready = icache_to_sram_r_ready; // @[Connect.scala 17:22]
  assign sram_i2_clock = clock;
  assign sram_i2_reset = reset;
  assign sram_i2_axi_ar_valid = EXU_i_lsu_axi_master_ar_valid; // @[Connect.scala 16:22]
  assign sram_i2_axi_ar_bits_addr = EXU_i_lsu_axi_master_ar_bits_addr; // @[Connect.scala 15:22]
  assign sram_i2_axi_r_ready = EXU_i_lsu_axi_master_r_ready; // @[Connect.scala 17:22]
  assign sram_i2_axi_aw_valid = EXU_i_lsu_axi_master_aw_valid; // @[Connect.scala 16:22]
  assign sram_i2_axi_aw_bits_addr = EXU_i_lsu_axi_master_aw_bits_addr; // @[Connect.scala 15:22]
  assign sram_i2_axi_w_valid = EXU_i_lsu_axi_master_w_valid; // @[Connect.scala 16:22]
  assign sram_i2_axi_w_bits_data = EXU_i_lsu_axi_master_w_bits_data; // @[Connect.scala 15:22]
  assign sram_i2_axi_w_bits_strb = EXU_i_lsu_axi_master_w_bits_strb; // @[Connect.scala 15:22]
  assign sram_i2_axi_b_ready = EXU_i_lsu_axi_master_b_ready; // @[Connect.scala 17:22]
  always @(posedge clock) begin
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_imm <= ISU_i_to_EXU_bits_imm; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_pc <= ISU_i_to_EXU_bits_pc; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_rdata1 <= ISU_i_to_EXU_bits_rdata1; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_rdata2 <= ISU_i_to_EXU_bits_rdata2; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_rd <= ISU_i_to_EXU_bits_rd; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen <= ISU_i_to_EXU_bits_ctrl_sig_reg_wen; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_fu_op <= ISU_i_to_EXU_bits_ctrl_sig_fu_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen <= ISU_i_to_EXU_bits_ctrl_sig_mem_wen; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak <= ISU_i_to_EXU_bits_ctrl_sig_is_ebreak; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_not_impl <= ISU_i_to_EXU_bits_ctrl_sig_not_impl; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_src1_op <= ISU_i_to_EXU_bits_ctrl_sig_src1_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_src2_op <= ISU_i_to_EXU_bits_ctrl_sig_src2_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_alu_op <= ISU_i_to_EXU_bits_ctrl_sig_alu_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op <= ISU_i_to_EXU_bits_ctrl_sig_lsu_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_bru_op <= ISU_i_to_EXU_bits_ctrl_sig_bru_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_csr_op <= ISU_i_to_EXU_bits_ctrl_sig_csr_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op <= ISU_i_to_EXU_bits_ctrl_sig_mdu_op; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_imm = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_rdata1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_rdata2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_rd = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_fu_op = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_not_impl = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_src1_op = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_src2_op = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_alu_op = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_bru_op = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_csr_op = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op = _RAND_16[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
