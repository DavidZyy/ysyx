
module memory (
    input      clk,
    input [] 
);
    
endmodule //memory
