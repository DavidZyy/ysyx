
`include "./include/defines.v"

module EX_MEM (
  
);
    
endmodule //EX_MEM
