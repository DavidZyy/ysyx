/* verilator lint_off DECLFILENAME */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off UNDRIVEN */
/* verilator lint_off UNOPTFLAT */
/* verilator lint_off WIDTHEXPAND */
module IDU(
  input         from_IFU_valid,
  input  [31:0] from_IFU_bits_inst,
  input  [31:0] from_IFU_bits_pc,
  output        to_ISU_valid,
  output [31:0] to_ISU_bits_imm,
  output [31:0] to_ISU_bits_pc,
  output [4:0]  to_ISU_bits_rs1,
  output [4:0]  to_ISU_bits_rs2,
  output [4:0]  to_ISU_bits_rd,
  output        to_ISU_bits_ctrl_sig_reg_wen,
  output [2:0]  to_ISU_bits_ctrl_sig_fu_op,
  output        to_ISU_bits_ctrl_sig_mem_wen,
  output        to_ISU_bits_ctrl_sig_is_ebreak,
  output        to_ISU_bits_ctrl_sig_not_impl,
  output [1:0]  to_ISU_bits_ctrl_sig_src1_op,
  output [1:0]  to_ISU_bits_ctrl_sig_src2_op,
  output [3:0]  to_ISU_bits_ctrl_sig_alu_op,
  output [3:0]  to_ISU_bits_ctrl_sig_lsu_op,
  output [3:0]  to_ISU_bits_ctrl_sig_bru_op,
  output [2:0]  to_ISU_bits_ctrl_sig_csr_op,
  output [3:0]  to_ISU_bits_ctrl_sig_mdu_op
);
  wire [19:0] _imm_i_T_2 = from_IFU_bits_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_i = {_imm_i_T_2,from_IFU_bits_inst[31:20]}; // @[Cat.scala 33:92]
  wire [31:0] imm_s = {_imm_i_T_2,from_IFU_bits_inst[31:25],from_IFU_bits_inst[11:7]}; // @[Cat.scala 33:92]
  wire [31:0] imm_b = {_imm_i_T_2,from_IFU_bits_inst[7],from_IFU_bits_inst[30:25],from_IFU_bits_inst[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] imm_u = {from_IFU_bits_inst[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [11:0] _imm_j_T_2 = from_IFU_bits_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 77:12]
  wire [32:0] imm_j = {_imm_j_T_2,from_IFU_bits_inst[31],from_IFU_bits_inst[19:12],from_IFU_bits_inst[20],
    from_IFU_bits_inst[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] decode_info_invInputs = ~from_IFU_bits_inst; // @[pla.scala 78:21]
  wire  decode_info_andMatrixInput_0 = from_IFU_bits_inst[0]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_1 = from_IFU_bits_inst[1]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_2 = decode_info_invInputs[2]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_3 = decode_info_invInputs[3]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_4 = decode_info_invInputs[4]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_5 = decode_info_invInputs[5]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_6 = decode_info_invInputs[6]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_7 = decode_info_invInputs[13]; // @[pla.scala 91:29]
  wire [7:0] _decode_info_T = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_1 = &_decode_info_T; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_6_1 = decode_info_invInputs[12]; // @[pla.scala 91:29]
  wire [7:0] _decode_info_T_2 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_3 = &_decode_info_T_2; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_7_2 = decode_info_invInputs[14]; // @[pla.scala 91:29]
  wire [7:0] _decode_info_T_4 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_5 = &_decode_info_T_4; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_6 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_7 = &_decode_info_T_6; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_8 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2,
    decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_9 = &_decode_info_T_8; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_10 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_6,decode_info_andMatrixInput_7
    ,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_11 = &_decode_info_T_10; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_4_6 = from_IFU_bits_inst[4]; // @[pla.scala 90:45]
  wire [7:0] _decode_info_T_12 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1}; // @[Cat.scala 33:92]
  wire  _decode_info_T_13 = &_decode_info_T_12; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_2_7 = from_IFU_bits_inst[2]; // @[pla.scala 90:45]
  wire [5:0] _decode_info_T_14 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_info_T_15 = &_decode_info_T_14; // @[pla.scala 98:74]
  wire [6:0] _decode_info_T_16 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_info_T_17 = &_decode_info_T_16; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_5_9 = from_IFU_bits_inst[5]; // @[pla.scala 90:45]
  wire [8:0] _decode_info_T_18 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_19 = &_decode_info_T_18; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_20 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_21 = &_decode_info_T_20; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_22 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_23 = &_decode_info_T_22; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_10 = decode_info_invInputs[25]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_11 = decode_info_invInputs[26]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_12 = decode_info_invInputs[27]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_13 = decode_info_invInputs[28]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_14 = decode_info_invInputs[29]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_15 = decode_info_invInputs[31]; // @[pla.scala 91:29]
  wire [7:0] decode_info_lo_12 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2,
    decode_info_andMatrixInput_10,decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,
    decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_24 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_12}; // @[Cat.scala 33:92]
  wire  _decode_info_T_25 = &_decode_info_T_24; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_11_1 = decode_info_invInputs[30]; // @[pla.scala 91:29]
  wire [5:0] decode_info_lo_13 = {decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,
    decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,
    decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [12:0] _decode_info_T_26 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_lo_13}; // @[Cat.scala 33:92]
  wire  _decode_info_T_27 = &_decode_info_T_26; // @[pla.scala 98:74]
  wire [6:0] decode_info_lo_14 = {decode_info_andMatrixInput_10,decode_info_andMatrixInput_11,
    decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,
    decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_T_28 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_lo_14}; // @[Cat.scala 33:92]
  wire  _decode_info_T_29 = &_decode_info_T_28; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_15 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_30 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_15}; // @[Cat.scala 33:92]
  wire  _decode_info_T_31 = &_decode_info_T_30; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_6_15 = from_IFU_bits_inst[6]; // @[pla.scala 90:45]
  wire [7:0] _decode_info_T_32 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_33 = &_decode_info_T_32; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_34 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_35 = &_decode_info_T_34; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_36 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_3
    ,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,
    decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_37 = &_decode_info_T_36; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_38 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_39 = &_decode_info_T_38; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_3_20 = from_IFU_bits_inst[3]; // @[pla.scala 90:45]
  wire [6:0] _decode_info_T_40 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2_7,decode_info_andMatrixInput_3_20,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15}; // @[Cat.scala 33:92]
  wire  _decode_info_T_41 = &_decode_info_T_40; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_7_18 = decode_info_invInputs[7]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_8_10 = decode_info_invInputs[8]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_9_5 = decode_info_invInputs[9]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_10_4 = decode_info_invInputs[10]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_11_4 = decode_info_invInputs[11]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_15_2 = decode_info_invInputs[15]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_16 = decode_info_invInputs[16]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_17 = decode_info_invInputs[17]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_18 = decode_info_invInputs[18]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_19 = decode_info_invInputs[19]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_20 = decode_info_invInputs[21]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_21 = decode_info_invInputs[22]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_22 = decode_info_invInputs[23]; // @[pla.scala 91:29]
  wire  decode_info_andMatrixInput_23 = decode_info_invInputs[24]; // @[pla.scala 91:29]
  wire [14:0] decode_info_lo_21 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,decode_info_andMatrixInput_20,
    decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_andMatrixInput_23,decode_info_lo_14}; // @[Cat.scala 33:92]
  wire [7:0] decode_info_hi_lo_20 = {decode_info_andMatrixInput_8_10,decode_info_andMatrixInput_9_5,
    decode_info_andMatrixInput_10_4,decode_info_andMatrixInput_11_4,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_15_2}; // @[Cat.scala 33:92]
  wire [30:0] _decode_info_T_42 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_21}; // @[Cat.scala 33:92]
  wire  _decode_info_T_43 = &_decode_info_T_42; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_20_1 = decode_info_invInputs[20]; // @[pla.scala 91:29]
  wire [7:0] decode_info_lo_lo_19 = {decode_info_andMatrixInput_23,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] decode_info_lo_22 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,decode_info_andMatrixInput_20_1,
    decode_info_andMatrixInput_20,decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_lo_lo_19}; // @[Cat.scala 33:92]
  wire [31:0] _decode_info_T_44 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_22}; // @[Cat.scala 33:92]
  wire  _decode_info_T_45 = &_decode_info_T_44; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_6_22 = from_IFU_bits_inst[12]; // @[pla.scala 90:45]
  wire [8:0] _decode_info_T_46 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_6,
    decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_47 = &_decode_info_T_46; // @[pla.scala 98:74]
  wire [6:0] decode_info_lo_24 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_11,
    decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,
    decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_T_48 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_24}; // @[Cat.scala 33:92]
  wire  _decode_info_T_49 = &_decode_info_T_48; // @[pla.scala 98:74]
  wire [14:0] _decode_info_T_50 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_24}; // @[Cat.scala 33:92]
  wire  _decode_info_T_51 = &_decode_info_T_50; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_52 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_53 = &_decode_info_T_52; // @[pla.scala 98:74]
  wire [15:0] _decode_info_T_54 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_15}; // @[Cat.scala 33:92]
  wire  _decode_info_T_55 = &_decode_info_T_54; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_56 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7}; // @[Cat.scala 33:92]
  wire  _decode_info_T_57 = &_decode_info_T_56; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_58 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,
    decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_59 = &_decode_info_T_58; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_60 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_61 = &_decode_info_T_60; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_8_20 = from_IFU_bits_inst[13]; // @[pla.scala 90:45]
  wire [9:0] _decode_info_T_62 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6
    ,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_63 = &_decode_info_T_62; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_64 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_8_20}; // @[Cat.scala 33:92]
  wire  _decode_info_T_65 = &_decode_info_T_64; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_66 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_67 = &_decode_info_T_66; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_68 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_20,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_69 = &_decode_info_T_68; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_35 = {decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_70 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_8_20,decode_info_lo_35}; // @[Cat.scala 33:92]
  wire  _decode_info_T_71 = &_decode_info_T_70; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_72 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_20,
    decode_info_andMatrixInput_7_2}; // @[Cat.scala 33:92]
  wire  _decode_info_T_73 = &_decode_info_T_72; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_74 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_8_20}; // @[Cat.scala 33:92]
  wire  _decode_info_T_75 = &_decode_info_T_74; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_38 = {decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_76 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_38}; // @[Cat.scala 33:92]
  wire  _decode_info_T_77 = &_decode_info_T_76; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_8_27 = from_IFU_bits_inst[14]; // @[pla.scala 90:45]
  wire [8:0] _decode_info_T_78 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6
    ,decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_79 = &_decode_info_T_78; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_80 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,decode_info_andMatrixInput_5,
    decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_81 = &_decode_info_T_80; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_41 = {decode_info_andMatrixInput_8_27,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_82 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_41}; // @[Cat.scala 33:92]
  wire  _decode_info_T_83 = &_decode_info_T_82; // @[pla.scala 98:74]
  wire [15:0] _decode_info_T_84 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_7,decode_info_lo_41}; // @[Cat.scala 33:92]
  wire  _decode_info_T_85 = &_decode_info_T_84; // @[pla.scala 98:74]
  wire [7:0] _decode_info_T_86 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_87 = &_decode_info_T_86; // @[pla.scala 98:74]
  wire [8:0] _decode_info_T_88 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_89 = &_decode_info_T_88; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_90 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5,decode_info_andMatrixInput_6
    ,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_91 = &_decode_info_T_90; // @[pla.scala 98:74]
  wire [6:0] decode_info_lo_46 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [14:0] _decode_info_T_92 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_46}; // @[Cat.scala 33:92]
  wire  _decode_info_T_93 = &_decode_info_T_92; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_47 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_94 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_47}; // @[Cat.scala 33:92]
  wire  _decode_info_T_95 = &_decode_info_T_94; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_48 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_10,decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,
    decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_96 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_48}; // @[Cat.scala 33:92]
  wire  _decode_info_T_97 = &_decode_info_T_96; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_98 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,decode_info_andMatrixInput_2
    ,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,decode_info_andMatrixInput_5_9,
    decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,decode_info_andMatrixInput_7,
    decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_99 = &_decode_info_T_98; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_100 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_101 = &_decode_info_T_100; // @[pla.scala 98:74]
  wire [9:0] _decode_info_T_102 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_8_27}; // @[Cat.scala 33:92]
  wire  _decode_info_T_103 = &_decode_info_T_102; // @[pla.scala 98:74]
  wire [15:0] decode_info_lo_52 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,from_IFU_bits_inst[20],decode_info_andMatrixInput_20,
    decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_lo_lo_19}; // @[Cat.scala 33:92]
  wire [31:0] _decode_info_T_104 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_52}; // @[Cat.scala 33:92]
  wire  _decode_info_T_105 = &_decode_info_T_104; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_7_50 = from_IFU_bits_inst[25]; // @[pla.scala 90:45]
  wire [6:0] decode_info_lo_53 = {decode_info_andMatrixInput_7_50,decode_info_andMatrixInput_11,
    decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,decode_info_andMatrixInput_14,
    decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_T_106 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_lo_53}; // @[Cat.scala 33:92]
  wire  _decode_info_T_107 = &_decode_info_T_106; // @[pla.scala 98:74]
  wire [14:0] _decode_info_T_108 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_53}; // @[Cat.scala 33:92]
  wire  _decode_info_T_109 = &_decode_info_T_108; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_55 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_110 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_55}; // @[Cat.scala 33:92]
  wire  _decode_info_T_111 = &_decode_info_T_110; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_56 = {decode_info_andMatrixInput_8_20,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_112 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_56}; // @[Cat.scala 33:92]
  wire  _decode_info_T_113 = &_decode_info_T_112; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_57 = {decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [16:0] _decode_info_T_114 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_8_20,decode_info_lo_57}; // @[Cat.scala 33:92]
  wire  _decode_info_T_115 = &_decode_info_T_114; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_58 = {decode_info_andMatrixInput_8_27,decode_info_andMatrixInput_7_50,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_116 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,decode_info_lo_58}; // @[Cat.scala 33:92]
  wire  _decode_info_T_117 = &_decode_info_T_116; // @[pla.scala 98:74]
  wire [15:0] _decode_info_T_118 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_7,decode_info_lo_58}; // @[Cat.scala 33:92]
  wire  _decode_info_T_119 = &_decode_info_T_118; // @[pla.scala 98:74]
  wire [16:0] _decode_info_T_120 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_8_20,decode_info_lo_58}; // @[Cat.scala 33:92]
  wire  _decode_info_T_121 = &_decode_info_T_120; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_21_3 = from_IFU_bits_inst[21]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_28_3 = from_IFU_bits_inst[28]; // @[pla.scala 90:45]
  wire  decode_info_andMatrixInput_29_3 = from_IFU_bits_inst[29]; // @[pla.scala 90:45]
  wire [7:0] decode_info_lo_lo_58 = {decode_info_andMatrixInput_23,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_28_3,
    decode_info_andMatrixInput_29_3,decode_info_andMatrixInput_11_1,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] decode_info_lo_61 = {decode_info_andMatrixInput_16,decode_info_andMatrixInput_17,
    decode_info_andMatrixInput_18,decode_info_andMatrixInput_19,decode_info_andMatrixInput_20_1,
    decode_info_andMatrixInput_21_3,decode_info_andMatrixInput_21,decode_info_andMatrixInput_22,decode_info_lo_lo_58}; // @[Cat.scala 33:92]
  wire [31:0] _decode_info_T_122 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6_15,decode_info_andMatrixInput_7_18,decode_info_hi_lo_20,
    decode_info_lo_61}; // @[Cat.scala 33:92]
  wire  _decode_info_T_123 = &_decode_info_T_122; // @[pla.scala 98:74]
  wire  decode_info_andMatrixInput_15_19 = from_IFU_bits_inst[30]; // @[pla.scala 90:45]
  wire [7:0] decode_info_lo_62 = {decode_info_andMatrixInput_7_2,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15_19,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [16:0] _decode_info_T_124 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_1,
    decode_info_andMatrixInput_7,decode_info_lo_62}; // @[Cat.scala 33:92]
  wire  _decode_info_T_125 = &_decode_info_T_124; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_63 = {decode_info_andMatrixInput_7,decode_info_andMatrixInput_8_27,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15_19,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [15:0] _decode_info_T_126 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,decode_info_lo_63}; // @[Cat.scala 33:92]
  wire  _decode_info_T_127 = &_decode_info_T_126; // @[pla.scala 98:74]
  wire [7:0] decode_info_lo_64 = {decode_info_andMatrixInput_8_27,decode_info_andMatrixInput_10,
    decode_info_andMatrixInput_11,decode_info_andMatrixInput_12,decode_info_andMatrixInput_13,
    decode_info_andMatrixInput_14,decode_info_andMatrixInput_15_19,decode_info_andMatrixInput_15}; // @[Cat.scala 33:92]
  wire [16:0] _decode_info_T_128 = {decode_info_andMatrixInput_0,decode_info_andMatrixInput_1,
    decode_info_andMatrixInput_2,decode_info_andMatrixInput_3,decode_info_andMatrixInput_4_6,
    decode_info_andMatrixInput_5_9,decode_info_andMatrixInput_6,decode_info_andMatrixInput_6_22,
    decode_info_andMatrixInput_7,decode_info_lo_64}; // @[Cat.scala 33:92]
  wire  _decode_info_T_129 = &_decode_info_T_128; // @[pla.scala 98:74]
  wire  _decode_info_orMatrixOutputs_T = |_decode_info_T_109; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_1 = {_decode_info_T_111,_decode_info_T_113}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_2 = |_decode_info_orMatrixOutputs_T_1; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_3 = {_decode_info_T_115,_decode_info_T_117,_decode_info_T_119}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_4 = |_decode_info_orMatrixOutputs_T_3; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_5 = |_decode_info_T_121; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_6 = {_decode_info_T_45,_decode_info_T_61}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_7 = |_decode_info_orMatrixOutputs_T_6; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_8 = {_decode_info_T_61,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_9 = |_decode_info_orMatrixOutputs_T_8; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_10 = |_decode_info_T_73; // @[pla.scala 114:39]
  wire [8:0] decode_info_orMatrixOutputs_lo = {_decode_info_T_43,_decode_info_T_49,_decode_info_T_59,_decode_info_T_65,
    _decode_info_T_73,_decode_info_T_87,_decode_info_T_93,_decode_info_T_97,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [17:0] _decode_info_orMatrixOutputs_T_11 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_11,
    _decode_info_T_15,_decode_info_T_25,_decode_info_T_27,_decode_info_T_37,_decode_info_T_41,
    decode_info_orMatrixOutputs_lo}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_12 = |_decode_info_orMatrixOutputs_T_11; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_13 = |_decode_info_T_105; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_14 = {_decode_info_T_19,_decode_info_T_23}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_15 = |_decode_info_orMatrixOutputs_T_14; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_1 = {_decode_info_T_41,_decode_info_T_49,_decode_info_T_61,_decode_info_T_65
    ,_decode_info_T_73,_decode_info_T_93,_decode_info_T_97}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_orMatrixOutputs_T_16 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_7,_decode_info_T_15,
    _decode_info_T_25,_decode_info_T_27,_decode_info_T_39,decode_info_orMatrixOutputs_lo_1}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_17 = |_decode_info_orMatrixOutputs_T_16; // @[pla.scala 114:39]
  wire [4:0] decode_info_orMatrixOutputs_lo_2 = {_decode_info_T_41,_decode_info_T_51,_decode_info_T_65,_decode_info_T_87
    ,_decode_info_T_93}; // @[Cat.scala 33:92]
  wire [10:0] _decode_info_orMatrixOutputs_T_18 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_15,
    _decode_info_T_21,_decode_info_T_37,decode_info_orMatrixOutputs_lo_2}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_19 = |_decode_info_orMatrixOutputs_T_18; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_3 = {_decode_info_T_37,_decode_info_T_41,_decode_info_T_49,_decode_info_T_65
    ,_decode_info_T_87,_decode_info_T_93,_decode_info_T_97}; // @[Cat.scala 33:92]
  wire [13:0] _decode_info_orMatrixOutputs_T_20 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_15,
    _decode_info_T_21,_decode_info_T_25,_decode_info_T_27,decode_info_orMatrixOutputs_lo_3}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_21 = |_decode_info_orMatrixOutputs_T_20; // @[pla.scala 114:39]
  wire [3:0] _decode_info_orMatrixOutputs_T_22 = {_decode_info_T_17,_decode_info_T_33,_decode_info_T_41,
    _decode_info_T_87}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_23 = |_decode_info_orMatrixOutputs_T_22; // @[pla.scala 114:39]
  wire [4:0] decode_info_orMatrixOutputs_lo_5 = {_decode_info_T_39,_decode_info_T_49,_decode_info_T_65,_decode_info_T_93
    ,_decode_info_T_97}; // @[Cat.scala 33:92]
  wire [10:0] _decode_info_orMatrixOutputs_T_24 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_11,
    _decode_info_T_25,_decode_info_T_27,decode_info_orMatrixOutputs_lo_5}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_25 = |_decode_info_orMatrixOutputs_T_24; // @[pla.scala 114:39]
  wire [5:0] decode_info_orMatrixOutputs_lo_6 = {_decode_info_T_41,_decode_info_T_75,_decode_info_T_77,_decode_info_T_85
    ,_decode_info_T_87,_decode_info_T_95}; // @[Cat.scala 33:92]
  wire [12:0] _decode_info_orMatrixOutputs_T_26 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_15,
    _decode_info_T_21,_decode_info_T_31,_decode_info_T_37,decode_info_orMatrixOutputs_lo_6}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_27 = |_decode_info_orMatrixOutputs_T_26; // @[pla.scala 114:39]
  wire [6:0] _decode_info_orMatrixOutputs_T_28 = {_decode_info_T_67,_decode_info_T_71,_decode_info_T_75,
    _decode_info_T_77,_decode_info_T_125,_decode_info_T_127,_decode_info_T_129}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_29 = |_decode_info_orMatrixOutputs_T_28; // @[pla.scala 114:39]
  wire [3:0] _decode_info_orMatrixOutputs_T_30 = {_decode_info_T_67,_decode_info_T_71,_decode_info_T_81,
    _decode_info_T_83}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_31 = |_decode_info_orMatrixOutputs_T_30; // @[pla.scala 114:39]
  wire [3:0] _decode_info_orMatrixOutputs_T_32 = {_decode_info_T_51,_decode_info_T_55,_decode_info_T_93,
    _decode_info_T_97}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_33 = |_decode_info_orMatrixOutputs_T_32; // @[pla.scala 114:39]
  wire [5:0] decode_info_orMatrixOutputs_lo_10 = {_decode_info_T_59,_decode_info_T_65,_decode_info_T_73,
    _decode_info_T_87,_decode_info_T_93,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [11:0] _decode_info_orMatrixOutputs_T_34 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_7,_decode_info_T_37,
    _decode_info_T_41,_decode_info_T_51,decode_info_orMatrixOutputs_lo_10}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_35 = |_decode_info_orMatrixOutputs_T_34; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_11 = {_decode_info_T_49,_decode_info_T_61,_decode_info_T_65,
    _decode_info_T_73,_decode_info_T_93,_decode_info_T_97,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [14:0] _decode_info_orMatrixOutputs_T_36 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_7,_decode_info_T_15,
    _decode_info_T_25,_decode_info_T_27,_decode_info_T_39,_decode_info_T_41,decode_info_orMatrixOutputs_lo_11}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_37 = |_decode_info_orMatrixOutputs_T_36; // @[pla.scala 114:39]
  wire [6:0] decode_info_orMatrixOutputs_lo_12 = {_decode_info_T_59,_decode_info_T_65,_decode_info_T_73,
    _decode_info_T_87,_decode_info_T_93,_decode_info_T_97,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire [14:0] _decode_info_orMatrixOutputs_T_38 = {_decode_info_T_1,_decode_info_T_3,_decode_info_T_5,_decode_info_T_11,
    _decode_info_T_25,_decode_info_T_27,_decode_info_T_37,_decode_info_T_49,decode_info_orMatrixOutputs_lo_12}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_39 = |_decode_info_orMatrixOutputs_T_38; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_40 = {_decode_info_T_35,_decode_info_T_41,_decode_info_T_89}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_41 = |_decode_info_orMatrixOutputs_T_40; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_42 = {_decode_info_T_37,_decode_info_T_99,_decode_info_T_101}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_43 = |_decode_info_orMatrixOutputs_T_42; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_44 = {_decode_info_T_57,_decode_info_T_89}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_45 = |_decode_info_orMatrixOutputs_T_44; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_46 = |_decode_info_T_103; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_47 = {_decode_info_T_9,_decode_info_T_53,_decode_info_T_91}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_48 = |_decode_info_orMatrixOutputs_T_47; // @[pla.scala 114:39]
  wire [2:0] _decode_info_orMatrixOutputs_T_49 = {_decode_info_T_23,_decode_info_T_47,_decode_info_T_63}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_50 = |_decode_info_orMatrixOutputs_T_49; // @[pla.scala 114:39]
  wire [1:0] _decode_info_orMatrixOutputs_T_51 = {_decode_info_T_23,_decode_info_T_79}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_52 = |_decode_info_orMatrixOutputs_T_51; // @[pla.scala 114:39]
  wire  _decode_info_orMatrixOutputs_T_53 = |_decode_info_T_69; // @[pla.scala 114:39]
  wire [14:0] _decode_info_orMatrixOutputs_T_54 = {_decode_info_T_13,_decode_info_T_15,_decode_info_T_25,
    _decode_info_T_29,_decode_info_T_37,_decode_info_T_41,_decode_info_T_43,_decode_info_T_51,
    decode_info_orMatrixOutputs_lo_12}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_55 = |_decode_info_orMatrixOutputs_T_54; // @[pla.scala 114:39]
  wire [4:0] _decode_info_orMatrixOutputs_T_56 = {_decode_info_T_33,_decode_info_T_37,_decode_info_T_41,
    _decode_info_T_87,_decode_info_T_107}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_57 = |_decode_info_orMatrixOutputs_T_56; // @[pla.scala 114:39]
  wire [6:0] _decode_info_orMatrixOutputs_T_58 = {_decode_info_T_1,_decode_info_T_5,_decode_info_T_11,_decode_info_T_43,
    _decode_info_T_61,_decode_info_T_73,_decode_info_T_123}; // @[Cat.scala 33:92]
  wire  _decode_info_orMatrixOutputs_T_59 = |_decode_info_orMatrixOutputs_T_58; // @[pla.scala 114:39]
  wire [7:0] decode_info_orMatrixOutputs_lo_lo_10 = {_decode_info_orMatrixOutputs_T_12,_decode_info_orMatrixOutputs_T_10
    ,_decode_info_orMatrixOutputs_T_9,_decode_info_orMatrixOutputs_T_7,_decode_info_orMatrixOutputs_T_5,
    _decode_info_orMatrixOutputs_T_4,_decode_info_orMatrixOutputs_T_2,_decode_info_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decode_info_orMatrixOutputs_hi_lo_12 = {_decode_info_orMatrixOutputs_T_43,_decode_info_orMatrixOutputs_T_41
    ,_decode_info_orMatrixOutputs_T_39,_decode_info_orMatrixOutputs_T_37,_decode_info_orMatrixOutputs_T_35,
    _decode_info_orMatrixOutputs_T_33,_decode_info_orMatrixOutputs_T_31,_decode_info_orMatrixOutputs_T_29}; // @[Cat.scala 33:92]
  wire [16:0] decode_info_orMatrixOutputs_hi_21 = {_decode_info_orMatrixOutputs_T_59,_decode_info_orMatrixOutputs_T_57,
    _decode_info_orMatrixOutputs_T_55,_decode_info_orMatrixOutputs_T_53,_decode_info_orMatrixOutputs_T_52,
    _decode_info_orMatrixOutputs_T_50,_decode_info_orMatrixOutputs_T_48,_decode_info_orMatrixOutputs_T_46,
    _decode_info_orMatrixOutputs_T_45,decode_info_orMatrixOutputs_hi_lo_12}; // @[Cat.scala 33:92]
  wire [32:0] decode_info_orMatrixOutputs = {decode_info_orMatrixOutputs_hi_21,_decode_info_orMatrixOutputs_T_27,
    _decode_info_orMatrixOutputs_T_25,_decode_info_orMatrixOutputs_T_23,_decode_info_orMatrixOutputs_T_21,
    _decode_info_orMatrixOutputs_T_19,_decode_info_orMatrixOutputs_T_17,_decode_info_orMatrixOutputs_T_15,
    _decode_info_orMatrixOutputs_T_13,decode_info_orMatrixOutputs_lo_lo_10}; // @[Cat.scala 33:92]
  wire  _decode_info_invMatrixOutputs_T_8 = ~decode_info_orMatrixOutputs[7]; // @[pla.scala 123:40]
  wire  _decode_info_invMatrixOutputs_T_22 = ~decode_info_orMatrixOutputs[20]; // @[pla.scala 123:40]
  wire  _decode_info_invMatrixOutputs_T_24 = ~decode_info_orMatrixOutputs[21]; // @[pla.scala 123:40]
  wire [7:0] decode_info_invMatrixOutputs_lo_lo = {_decode_info_invMatrixOutputs_T_8,decode_info_orMatrixOutputs[6],
    decode_info_orMatrixOutputs[5],decode_info_orMatrixOutputs[4],decode_info_orMatrixOutputs[3],
    decode_info_orMatrixOutputs[2],decode_info_orMatrixOutputs[1],decode_info_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] decode_info_invMatrixOutputs_hi_lo = {decode_info_orMatrixOutputs[23],decode_info_orMatrixOutputs[22],
    _decode_info_invMatrixOutputs_T_24,_decode_info_invMatrixOutputs_T_22,decode_info_orMatrixOutputs[19],
    decode_info_orMatrixOutputs[18],decode_info_orMatrixOutputs[17],decode_info_orMatrixOutputs[16]}; // @[Cat.scala 33:92]
  wire [16:0] decode_info_invMatrixOutputs_hi = {decode_info_orMatrixOutputs[32],decode_info_orMatrixOutputs[31],
    decode_info_orMatrixOutputs[30],decode_info_orMatrixOutputs[29],decode_info_orMatrixOutputs[28],
    decode_info_orMatrixOutputs[27],decode_info_orMatrixOutputs[26],decode_info_orMatrixOutputs[25],
    decode_info_orMatrixOutputs[24],decode_info_invMatrixOutputs_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] decode_info_invMatrixOutputs = {decode_info_invMatrixOutputs_hi,decode_info_orMatrixOutputs[15],
    decode_info_orMatrixOutputs[14],decode_info_orMatrixOutputs[13],decode_info_orMatrixOutputs[12],
    decode_info_orMatrixOutputs[11],decode_info_orMatrixOutputs[10],decode_info_orMatrixOutputs[9],
    decode_info_orMatrixOutputs[8],decode_info_invMatrixOutputs_lo_lo}; // @[Cat.scala 33:92]
  wire [2:0] inst_type = decode_info_invMatrixOutputs[21:19]; // @[IDU.scala 111:36]
  wire [31:0] _to_ISU_bits_imm_T_1 = 3'h1 == inst_type ? imm_i : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_imm_T_3 = 3'h2 == inst_type ? imm_s : _to_ISU_bits_imm_T_1; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_imm_T_5 = 3'h3 == inst_type ? imm_b : _to_ISU_bits_imm_T_3; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_imm_T_7 = 3'h4 == inst_type ? imm_u : _to_ISU_bits_imm_T_5; // @[Mux.scala 81:58]
  wire [32:0] _to_ISU_bits_imm_T_9 = 3'h5 == inst_type ? imm_j : {{1'd0}, _to_ISU_bits_imm_T_7}; // @[Mux.scala 81:58]
  assign to_ISU_valid = from_IFU_valid; // @[IDU.scala 17:20]
  assign to_ISU_bits_imm = _to_ISU_bits_imm_T_9[31:0]; // @[IDU.scala 112:21]
  assign to_ISU_bits_pc = from_IFU_bits_pc; // @[IDU.scala 122:21]
  assign to_ISU_bits_rs1 = from_IFU_bits_inst[19:15]; // @[IDU.scala 119:42]
  assign to_ISU_bits_rs2 = from_IFU_bits_inst[24:20]; // @[IDU.scala 120:42]
  assign to_ISU_bits_rd = from_IFU_bits_inst[11:7]; // @[IDU.scala 121:42]
  assign to_ISU_bits_ctrl_sig_reg_wen = decode_info_invMatrixOutputs[10]; // @[IDU.scala 130:50]
  assign to_ISU_bits_ctrl_sig_fu_op = decode_info_invMatrixOutputs[32:30]; // @[IDU.scala 136:50]
  assign to_ISU_bits_ctrl_sig_mem_wen = decode_info_invMatrixOutputs[9]; // @[IDU.scala 129:50]
  assign to_ISU_bits_ctrl_sig_is_ebreak = decode_info_invMatrixOutputs[8]; // @[IDU.scala 128:50]
  assign to_ISU_bits_ctrl_sig_not_impl = decode_info_invMatrixOutputs[7]; // @[IDU.scala 127:50]
  assign to_ISU_bits_ctrl_sig_src1_op = decode_info_invMatrixOutputs[14:13]; // @[IDU.scala 132:50]
  assign to_ISU_bits_ctrl_sig_src2_op = decode_info_invMatrixOutputs[12:11]; // @[IDU.scala 131:50]
  assign to_ISU_bits_ctrl_sig_alu_op = decode_info_invMatrixOutputs[18:15]; // @[IDU.scala 133:50]
  assign to_ISU_bits_ctrl_sig_lsu_op = decode_info_invMatrixOutputs[29:26]; // @[IDU.scala 135:50]
  assign to_ISU_bits_ctrl_sig_bru_op = decode_info_invMatrixOutputs[25:22]; // @[IDU.scala 134:50]
  assign to_ISU_bits_ctrl_sig_csr_op = decode_info_invMatrixOutputs[6:4]; // @[IDU.scala 126:50]
  assign to_ISU_bits_ctrl_sig_mdu_op = decode_info_invMatrixOutputs[3:0]; // @[IDU.scala 125:50]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_in_rs1,
  input  [4:0]  io_in_rs2,
  input  [4:0]  io_in_rd,
  input  [31:0] io_in_wdata,
  input         io_in_reg_wen,
  output [31:0] io_out_rdata1,
  output [31:0] io_out_rdata2
);
  wire  regfile_clock; // @[regfile.scala 48:25]
  wire  regfile_reset; // @[regfile.scala 48:25]
  wire [4:0] regfile_rs1; // @[regfile.scala 48:25]
  wire [4:0] regfile_rs2; // @[regfile.scala 48:25]
  wire [4:0] regfile_rd; // @[regfile.scala 48:25]
  wire [31:0] regfile_wdata; // @[regfile.scala 48:25]
  wire  regfile_reg_wen; // @[regfile.scala 48:25]
  wire [31:0] regfile_rdata1; // @[regfile.scala 48:25]
  wire [31:0] regfile_rdata2; // @[regfile.scala 48:25]
  RegisterFileBB regfile ( // @[regfile.scala 48:25]
    .clock(regfile_clock),
    .reset(regfile_reset),
    .rs1(regfile_rs1),
    .rs2(regfile_rs2),
    .rd(regfile_rd),
    .wdata(regfile_wdata),
    .reg_wen(regfile_reg_wen),
    .rdata1(regfile_rdata1),
    .rdata2(regfile_rdata2)
  );
  assign io_out_rdata1 = regfile_rdata1; // @[regfile.scala 58:19]
  assign io_out_rdata2 = regfile_rdata2; // @[regfile.scala 59:19]
  assign regfile_clock = clock; // @[regfile.scala 50:24]
  assign regfile_reset = reset; // @[regfile.scala 51:24]
  assign regfile_rs1 = io_in_rs1; // @[regfile.scala 52:24]
  assign regfile_rs2 = io_in_rs2; // @[regfile.scala 53:24]
  assign regfile_rd = io_in_rd; // @[regfile.scala 54:24]
  assign regfile_wdata = io_in_wdata; // @[regfile.scala 55:24]
  assign regfile_reg_wen = io_in_reg_wen; // @[regfile.scala 56:24]
endmodule
module ISU(
  input         clock,
  input         reset,
  input         from_IDU_valid,
  input  [31:0] from_IDU_bits_imm,
  input  [31:0] from_IDU_bits_pc,
  input  [4:0]  from_IDU_bits_rs1,
  input  [4:0]  from_IDU_bits_rs2,
  input  [4:0]  from_IDU_bits_rd,
  input         from_IDU_bits_ctrl_sig_reg_wen,
  input  [2:0]  from_IDU_bits_ctrl_sig_fu_op,
  input         from_IDU_bits_ctrl_sig_mem_wen,
  input         from_IDU_bits_ctrl_sig_is_ebreak,
  input         from_IDU_bits_ctrl_sig_not_impl,
  input  [1:0]  from_IDU_bits_ctrl_sig_src1_op,
  input  [1:0]  from_IDU_bits_ctrl_sig_src2_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_alu_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_lsu_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_bru_op,
  input  [2:0]  from_IDU_bits_ctrl_sig_csr_op,
  input  [3:0]  from_IDU_bits_ctrl_sig_mdu_op,
  input         from_WBU_bits_reg_wen,
  input  [31:0] from_WBU_bits_wdata,
  input  [4:0]  from_WBU_bits_rd,
  output        to_EXU_valid,
  output [31:0] to_EXU_bits_imm,
  output [31:0] to_EXU_bits_pc,
  output [31:0] to_EXU_bits_rdata1,
  output [31:0] to_EXU_bits_rdata2,
  output [4:0]  to_EXU_bits_rd,
  output        to_EXU_bits_ctrl_sig_reg_wen,
  output [2:0]  to_EXU_bits_ctrl_sig_fu_op,
  output        to_EXU_bits_ctrl_sig_mem_wen,
  output        to_EXU_bits_ctrl_sig_is_ebreak,
  output        to_EXU_bits_ctrl_sig_not_impl,
  output [1:0]  to_EXU_bits_ctrl_sig_src1_op,
  output [1:0]  to_EXU_bits_ctrl_sig_src2_op,
  output [3:0]  to_EXU_bits_ctrl_sig_alu_op,
  output [3:0]  to_EXU_bits_ctrl_sig_lsu_op,
  output [3:0]  to_EXU_bits_ctrl_sig_bru_op,
  output [2:0]  to_EXU_bits_ctrl_sig_csr_op,
  output [3:0]  to_EXU_bits_ctrl_sig_mdu_op
);
  wire  RegFile_i_clock; // @[ISU.scala 20:37]
  wire  RegFile_i_reset; // @[ISU.scala 20:37]
  wire [4:0] RegFile_i_io_in_rs1; // @[ISU.scala 20:37]
  wire [4:0] RegFile_i_io_in_rs2; // @[ISU.scala 20:37]
  wire [4:0] RegFile_i_io_in_rd; // @[ISU.scala 20:37]
  wire [31:0] RegFile_i_io_in_wdata; // @[ISU.scala 20:37]
  wire  RegFile_i_io_in_reg_wen; // @[ISU.scala 20:37]
  wire [31:0] RegFile_i_io_out_rdata1; // @[ISU.scala 20:37]
  wire [31:0] RegFile_i_io_out_rdata2; // @[ISU.scala 20:37]
  RegFile RegFile_i ( // @[ISU.scala 20:37]
    .clock(RegFile_i_clock),
    .reset(RegFile_i_reset),
    .io_in_rs1(RegFile_i_io_in_rs1),
    .io_in_rs2(RegFile_i_io_in_rs2),
    .io_in_rd(RegFile_i_io_in_rd),
    .io_in_wdata(RegFile_i_io_in_wdata),
    .io_in_reg_wen(RegFile_i_io_in_reg_wen),
    .io_out_rdata1(RegFile_i_io_out_rdata1),
    .io_out_rdata2(RegFile_i_io_out_rdata2)
  );
  assign to_EXU_valid = from_IDU_valid; // @[ISU.scala 18:20]
  assign to_EXU_bits_imm = from_IDU_bits_imm; // @[ISU.scala 33:26]
  assign to_EXU_bits_pc = from_IDU_bits_pc; // @[ISU.scala 34:26]
  assign to_EXU_bits_rdata1 = RegFile_i_io_out_rdata1; // @[ISU.scala 36:26]
  assign to_EXU_bits_rdata2 = RegFile_i_io_out_rdata2; // @[ISU.scala 37:26]
  assign to_EXU_bits_rd = from_IDU_bits_rd; // @[ISU.scala 35:26]
  assign to_EXU_bits_ctrl_sig_reg_wen = from_IDU_bits_ctrl_sig_reg_wen; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_fu_op = from_IDU_bits_ctrl_sig_fu_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_mem_wen = from_IDU_bits_ctrl_sig_mem_wen; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_is_ebreak = from_IDU_bits_ctrl_sig_is_ebreak; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_not_impl = from_IDU_bits_ctrl_sig_not_impl; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_src1_op = from_IDU_bits_ctrl_sig_src1_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_src2_op = from_IDU_bits_ctrl_sig_src2_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_alu_op = from_IDU_bits_ctrl_sig_alu_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_lsu_op = from_IDU_bits_ctrl_sig_lsu_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_bru_op = from_IDU_bits_ctrl_sig_bru_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_csr_op = from_IDU_bits_ctrl_sig_csr_op; // @[ISU.scala 32:26]
  assign to_EXU_bits_ctrl_sig_mdu_op = from_IDU_bits_ctrl_sig_mdu_op; // @[ISU.scala 32:26]
  assign RegFile_i_clock = clock;
  assign RegFile_i_reset = reset;
  assign RegFile_i_io_in_rs1 = from_IDU_bits_rs1; // @[ISU.scala 24:29]
  assign RegFile_i_io_in_rs2 = from_IDU_bits_rs2; // @[ISU.scala 25:29]
  assign RegFile_i_io_in_rd = from_WBU_bits_rd; // @[ISU.scala 23:29]
  assign RegFile_i_io_in_wdata = from_WBU_bits_wdata; // @[ISU.scala 29:29]
  assign RegFile_i_io_in_reg_wen = from_WBU_bits_reg_wen; // @[ISU.scala 28:29]
endmodule
module Alu(
  input  [31:0] io_in_src1,
  input  [31:0] io_in_src2,
  input  [3:0]  io_in_op,
  output [31:0] io_out_result
);
  wire [4:0] shamt = io_in_src2[4:0]; // @[alu.scala 31:25]
  wire [31:0] _io_out_result_T_1 = io_in_src1 + io_in_src2; // @[alu.scala 36:42]
  wire [31:0] _io_out_result_T_3 = io_in_src1 - io_in_src2; // @[alu.scala 37:42]
  wire [31:0] _io_out_result_T_4 = io_in_src1 & io_in_src2; // @[alu.scala 38:42]
  wire [31:0] _io_out_result_T_5 = io_in_src1 | io_in_src2; // @[alu.scala 39:42]
  wire [31:0] _io_out_result_T_6 = io_in_src1 ^ io_in_src2; // @[alu.scala 40:42]
  wire  _io_out_result_T_9 = $signed(io_in_src1) < $signed(io_in_src2); // @[alu.scala 41:49]
  wire  _io_out_result_T_10 = io_in_src1 < io_in_src2; // @[alu.scala 42:42]
  wire [62:0] _GEN_0 = {{31'd0}, io_in_src1}; // @[alu.scala 43:42]
  wire [62:0] _io_out_result_T_11 = _GEN_0 << shamt; // @[alu.scala 43:42]
  wire [31:0] _io_out_result_T_12 = io_in_src1 >> shamt; // @[alu.scala 44:42]
  wire [31:0] _io_out_result_T_15 = $signed(io_in_src1) >>> shamt; // @[alu.scala 45:59]
  wire [31:0] _io_out_result_T_19 = 4'h1 == io_in_op ? _io_out_result_T_1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_21 = 4'h2 == io_in_op ? _io_out_result_T_3 : _io_out_result_T_19; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_23 = 4'h3 == io_in_op ? _io_out_result_T_4 : _io_out_result_T_21; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_25 = 4'h4 == io_in_op ? _io_out_result_T_5 : _io_out_result_T_23; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_27 = 4'h5 == io_in_op ? _io_out_result_T_6 : _io_out_result_T_25; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_29 = 4'h6 == io_in_op ? {{31'd0}, _io_out_result_T_9} : _io_out_result_T_27; // @[Mux.scala 81:58]
  wire [31:0] _io_out_result_T_31 = 4'h7 == io_in_op ? {{31'd0}, _io_out_result_T_10} : _io_out_result_T_29; // @[Mux.scala 81:58]
  wire [62:0] _io_out_result_T_33 = 4'h8 == io_in_op ? _io_out_result_T_11 : {{31'd0}, _io_out_result_T_31}; // @[Mux.scala 81:58]
  wire [62:0] _io_out_result_T_35 = 4'h9 == io_in_op ? {{31'd0}, _io_out_result_T_12} : _io_out_result_T_33; // @[Mux.scala 81:58]
  wire [62:0] _io_out_result_T_37 = 4'ha == io_in_op ? {{31'd0}, _io_out_result_T_15} : _io_out_result_T_35; // @[Mux.scala 81:58]
  assign io_out_result = _io_out_result_T_37[31:0]; // @[alu.scala 33:21]
endmodule
module Mdu(
  input  [31:0] io_in_src1,
  input  [31:0] io_in_src2,
  input  [3:0]  io_in_op,
  output [31:0] io_out_result
);
  wire [63:0] _io_out_result_T = io_in_src1 * io_in_src2; // @[mdu.scala 36:44]
  wire [63:0] _io_out_result_T_3 = $signed(io_in_src1) * $signed(io_in_src2); // @[mdu.scala 37:52]
  wire [31:0] _io_out_result_T_5 = _io_out_result_T_3[63:32]; // @[mdu.scala 37:86]
  wire [32:0] _io_out_result_T_7 = {1'b0,$signed(io_in_src2)}; // @[mdu.scala 38:52]
  wire [64:0] _io_out_result_T_8 = $signed(io_in_src1) * $signed(_io_out_result_T_7); // @[mdu.scala 38:52]
  wire [63:0] _io_out_result_T_10 = _io_out_result_T_8[63:0]; // @[mdu.scala 38:52]
  wire [31:0] _io_out_result_T_12 = _io_out_result_T_10[63:32]; // @[mdu.scala 38:79]
  wire [32:0] _io_out_result_T_18 = $signed(io_in_src1) / $signed(io_in_src2); // @[mdu.scala 40:70]
  wire [31:0] _io_out_result_T_19 = io_in_src1 / io_in_src2; // @[mdu.scala 41:44]
  wire [31:0] _io_out_result_T_23 = $signed(io_in_src1) % $signed(io_in_src2); // @[mdu.scala 42:70]
  wire [31:0] _io_out_result_T_24 = io_in_src1 % io_in_src2; // @[mdu.scala 43:44]
  wire [63:0] _io_out_result_T_28 = 4'h1 == io_in_op ? _io_out_result_T : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_30 = 4'h2 == io_in_op ? {{32'd0}, _io_out_result_T_5} : _io_out_result_T_28; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_32 = 4'h3 == io_in_op ? {{32'd0}, _io_out_result_T_12} : _io_out_result_T_30; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_34 = 4'h4 == io_in_op ? {{32'd0}, _io_out_result_T[63:32]} : _io_out_result_T_32; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_36 = 4'h5 == io_in_op ? {{31'd0}, _io_out_result_T_18} : _io_out_result_T_34; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_38 = 4'h6 == io_in_op ? {{32'd0}, _io_out_result_T_19} : _io_out_result_T_36; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_40 = 4'h7 == io_in_op ? {{32'd0}, _io_out_result_T_23} : _io_out_result_T_38; // @[Mux.scala 81:58]
  wire [63:0] _io_out_result_T_42 = 4'h8 == io_in_op ? {{32'd0}, _io_out_result_T_24} : _io_out_result_T_40; // @[Mux.scala 81:58]
  assign io_out_result = _io_out_result_T_42[31:0]; // @[mdu.scala 33:21]
endmodule
module Bru(
  input  [31:0] io_in_src1,
  input  [31:0] io_in_src2,
  input  [3:0]  io_in_op,
  output        io_out_ctrl_br
);
  wire  _io_out_ctrl_br_T = io_in_src1 == io_in_src2; // @[bru.scala 35:44]
  wire  _io_out_ctrl_br_T_1 = io_in_src1 != io_in_src2; // @[bru.scala 36:44]
  wire  _io_out_ctrl_br_T_4 = $signed(io_in_src1) < $signed(io_in_src2); // @[bru.scala 37:51]
  wire  _io_out_ctrl_br_T_7 = $signed(io_in_src1) >= $signed(io_in_src2); // @[bru.scala 38:51]
  wire  _io_out_ctrl_br_T_8 = io_in_src1 < io_in_src2; // @[bru.scala 39:51]
  wire  _io_out_ctrl_br_T_9 = io_in_src1 >= io_in_src2; // @[bru.scala 40:51]
  wire  _io_out_ctrl_br_T_15 = 4'h3 == io_in_op ? _io_out_ctrl_br_T : 4'h2 == io_in_op | 4'h1 == io_in_op; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_17 = 4'h4 == io_in_op ? _io_out_ctrl_br_T_1 : _io_out_ctrl_br_T_15; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_19 = 4'h5 == io_in_op ? _io_out_ctrl_br_T_4 : _io_out_ctrl_br_T_17; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_21 = 4'h6 == io_in_op ? _io_out_ctrl_br_T_7 : _io_out_ctrl_br_T_19; // @[Mux.scala 81:58]
  wire  _io_out_ctrl_br_T_23 = 4'h7 == io_in_op ? _io_out_ctrl_br_T_8 : _io_out_ctrl_br_T_21; // @[Mux.scala 81:58]
  assign io_out_ctrl_br = 4'h8 == io_in_op ? _io_out_ctrl_br_T_9 : _io_out_ctrl_br_T_23; // @[Mux.scala 81:58]
endmodule
module Lsu(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_mem_wen,
  input  [31:0] io_in_addr,
  input  [31:0] io_in_wdata,
  input  [3:0]  io_in_op,
  output [31:0] io_out_rdata,
  output        io_out_end,
  output        io_out_idle,
  input         axi_ar_ready,
  output        axi_ar_valid,
  output [31:0] axi_ar_bits_addr,
  output        axi_r_ready,
  input         axi_r_valid,
  input  [31:0] axi_r_bits_data,
  input         axi_aw_ready,
  output        axi_aw_valid,
  output [31:0] axi_aw_bits_addr,
  input         axi_w_ready,
  output        axi_w_valid,
  output [31:0] axi_w_bits_data,
  output [3:0]  axi_w_bits_strb,
  output        axi_b_ready,
  input         axi_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[lsu.scala 35:24]
  wire  _state_T = axi_ar_ready & axi_ar_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_2 = axi_r_ready & axi_r_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_3 = _state_T_2 ? 3'h5 : 3'h2; // @[lsu.scala 53:25]
  wire  _state_T_4 = axi_aw_ready & axi_aw_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_5 = axi_w_ready & axi_w_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_7 = _state_T_4 & _state_T_5 ? 3'h4 : 3'h3; // @[lsu.scala 58:25]
  wire  _state_T_8 = axi_b_ready & axi_b_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_9 = _state_T_8 ? 3'h5 : 3'h4; // @[lsu.scala 61:25]
  wire [2:0] _GEN_2 = 3'h5 == state ? 3'h0 : state; // @[lsu.scala 36:20 64:19 35:24]
  wire [2:0] _GEN_3 = 3'h4 == state ? _state_T_9 : _GEN_2; // @[lsu.scala 36:20 61:19]
  wire [2:0] _GEN_4 = 3'h3 == state ? _state_T_7 : _GEN_3; // @[lsu.scala 36:20 58:19]
  wire [1:0] addr_low_2 = io_in_addr[1:0]; // @[lsu.scala 71:31]
  wire [23:0] _lb_rdata_T_2 = axi_r_bits_data[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_4 = {_lb_rdata_T_2,axi_r_bits_data[7:0]}; // @[Cat.scala 33:92]
  wire [23:0] _lb_rdata_T_7 = axi_r_bits_data[15] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_9 = {_lb_rdata_T_7,axi_r_bits_data[15:8]}; // @[Cat.scala 33:92]
  wire [23:0] _lb_rdata_T_12 = axi_r_bits_data[23] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_14 = {_lb_rdata_T_12,axi_r_bits_data[23:16]}; // @[Cat.scala 33:92]
  wire [23:0] _lb_rdata_T_17 = axi_r_bits_data[31] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lb_rdata_T_19 = {_lb_rdata_T_17,axi_r_bits_data[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _lb_rdata_T_21 = 2'h1 == addr_low_2 ? _lb_rdata_T_9 : _lb_rdata_T_4; // @[Mux.scala 81:58]
  wire [31:0] _lb_rdata_T_23 = 2'h2 == addr_low_2 ? _lb_rdata_T_14 : _lb_rdata_T_21; // @[Mux.scala 81:58]
  wire [31:0] lb_rdata = 2'h3 == addr_low_2 ? _lb_rdata_T_19 : _lb_rdata_T_23; // @[Mux.scala 81:58]
  wire [31:0] _lbu_rdata_T_2 = {24'h0,axi_r_bits_data[7:0]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_5 = {24'h0,axi_r_bits_data[15:8]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_8 = {24'h0,axi_r_bits_data[23:16]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_11 = {24'h0,axi_r_bits_data[31:24]}; // @[Cat.scala 33:92]
  wire [31:0] _lbu_rdata_T_13 = 2'h1 == addr_low_2 ? _lbu_rdata_T_5 : _lbu_rdata_T_2; // @[Mux.scala 81:58]
  wire [31:0] _lbu_rdata_T_15 = 2'h2 == addr_low_2 ? _lbu_rdata_T_8 : _lbu_rdata_T_13; // @[Mux.scala 81:58]
  wire [31:0] lbu_rdata = 2'h3 == addr_low_2 ? _lbu_rdata_T_11 : _lbu_rdata_T_15; // @[Mux.scala 81:58]
  wire [15:0] _lh_rdata_T_2 = axi_r_bits_data[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lh_rdata_T_4 = {_lh_rdata_T_2,axi_r_bits_data[15:0]}; // @[Cat.scala 33:92]
  wire [15:0] _lh_rdata_T_7 = axi_r_bits_data[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _lh_rdata_T_9 = {_lh_rdata_T_7,axi_r_bits_data[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _lh_rdata_T_11 = 2'h0 == addr_low_2 ? _lh_rdata_T_4 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] lh_rdata = 2'h2 == addr_low_2 ? _lh_rdata_T_9 : _lh_rdata_T_11; // @[Mux.scala 81:58]
  wire [31:0] _lhu_rdata_T_2 = {16'h0,axi_r_bits_data[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _lhu_rdata_T_5 = {16'h0,axi_r_bits_data[31:16]}; // @[Cat.scala 33:92]
  wire [31:0] _lhu_rdata_T_7 = 2'h0 == addr_low_2 ? _lhu_rdata_T_2 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] lhu_rdata = 2'h2 == addr_low_2 ? _lhu_rdata_T_5 : _lhu_rdata_T_7; // @[Mux.scala 81:58]
  wire [1:0] _sb_wmask_T_1 = 2'h1 == addr_low_2 ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [2:0] _sb_wmask_T_3 = 2'h2 == addr_low_2 ? 3'h4 : {{1'd0}, _sb_wmask_T_1}; // @[Mux.scala 81:58]
  wire [3:0] sb_wmask = 2'h3 == addr_low_2 ? 4'h8 : {{1'd0}, _sb_wmask_T_3}; // @[Mux.scala 81:58]
  wire [1:0] _sh_wmask_T_1 = 2'h0 == addr_low_2 ? 2'h3 : 2'h0; // @[Mux.scala 81:58]
  wire [3:0] sh_wmask = 2'h2 == addr_low_2 ? 4'hc : {{2'd0}, _sh_wmask_T_1}; // @[Mux.scala 81:58]
  wire [3:0] _wmask_T_1 = 4'h6 == io_in_op ? sb_wmask : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _wmask_T_3 = 4'h7 == io_in_op ? sh_wmask : _wmask_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_3 = 4'h1 == io_in_op ? lb_rdata : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_5 = 4'h4 == io_in_op ? lbu_rdata : _io_out_rdata_T_3; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_7 = 4'h2 == io_in_op ? lh_rdata : _io_out_rdata_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_out_rdata_T_9 = 4'h5 == io_in_op ? lhu_rdata : _io_out_rdata_T_7; // @[Mux.scala 81:58]
  assign io_out_rdata = 4'h3 == io_in_op ? axi_r_bits_data : _io_out_rdata_T_9; // @[Mux.scala 81:58]
  assign io_out_end = 3'h5 == state; // @[Mux.scala 81:61]
  assign io_out_idle = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_ar_valid = 3'h1 == state; // @[Mux.scala 81:61]
  assign axi_ar_bits_addr = io_in_addr; // @[lsu.scala 148:22]
  assign axi_r_ready = 3'h2 == state; // @[Mux.scala 81:61]
  assign axi_aw_valid = 3'h3 == state; // @[Mux.scala 81:61]
  assign axi_aw_bits_addr = io_in_addr; // @[lsu.scala 151:22]
  assign axi_w_valid = 3'h3 == state; // @[Mux.scala 81:61]
  assign axi_w_bits_data = io_in_wdata; // @[lsu.scala 153:22]
  assign axi_w_bits_strb = 4'h8 == io_in_op ? 4'hf : _wmask_T_3; // @[Mux.scala 81:58]
  assign axi_b_ready = 3'h4 == state; // @[Mux.scala 81:61]
  always @(posedge clock) begin
    if (reset) begin // @[lsu.scala 35:24]
      state <= 3'h0; // @[lsu.scala 35:24]
    end else if (3'h0 == state) begin // @[lsu.scala 36:20]
      if (io_in_valid) begin // @[lsu.scala 38:32]
        if (io_in_mem_wen) begin // @[lsu.scala 39:38]
          state <= 3'h3; // @[lsu.scala 40:27]
        end else begin
          state <= 3'h1; // @[lsu.scala 42:27]
        end
      end else begin
        state <= 3'h0; // @[lsu.scala 45:23]
      end
    end else if (3'h1 == state) begin // @[lsu.scala 36:20]
      if (_state_T) begin // @[lsu.scala 50:25]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[lsu.scala 36:20]
      state <= _state_T_3; // @[lsu.scala 53:19]
    end else begin
      state <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csr(
  input         clock,
  input         reset,
  input  [2:0]  io_in_op,
  input  [31:0] io_in_cur_pc,
  input  [31:0] io_in_csr_id,
  input  [31:0] io_in_wdata,
  output        io_out_csr_br,
  output [31:0] io_out_csr_addr,
  output [31:0] io_out_r_csr,
  output [31:0] io_out_difftest_mcause,
  output [31:0] io_out_difftest_mepc,
  output [31:0] io_out_difftest_mstatus,
  output [31:0] io_out_difftest_mtvec
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_mepc; // @[csr.scala 32:28]
  reg [31:0] reg_mcause; // @[csr.scala 33:28]
  reg [31:0] reg_mstatus; // @[csr.scala 34:28]
  reg [31:0] reg_mtvec; // @[csr.scala 35:28]
  wire [31:0] _reg_mcause_csrrs_T = io_in_wdata | reg_mcause; // @[csr.scala 51:32]
  wire [31:0] _reg_mepc_csrrs_T = io_in_wdata | reg_mepc; // @[csr.scala 63:30]
  wire [31:0] _reg_mstatus_csrrs_T = io_in_wdata | reg_mstatus; // @[csr.scala 75:33]
  wire [31:0] _reg_mstatus_T_5 = {reg_mstatus[31:13],2'h3,reg_mstatus[10:8],reg_mstatus[3],reg_mstatus[6:4],1'h0,
    reg_mstatus[2:0]}; // @[Cat.scala 33:92]
  wire [30:0] _reg_mstatus_T_11 = {reg_mstatus[31:13],1'h0,reg_mstatus[10:8],1'h1,reg_mstatus[6:4],reg_mstatus[7],
    reg_mstatus[2:0]}; // @[Cat.scala 33:92]
  wire [31:0] _reg_mstatus_T_13 = 3'h1 == io_in_op ? _reg_mstatus_T_5 : reg_mstatus; // @[Mux.scala 81:58]
  wire [31:0] _reg_mtvec_csrrs_T = io_in_wdata | reg_mtvec; // @[csr.scala 100:31]
  wire [31:0] _io_out_csr_addr_T_1 = 3'h1 == io_in_op ? reg_mtvec : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_r_csr_T_1 = 32'h305 == io_in_csr_id ? reg_mtvec : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_out_r_csr_T_3 = 32'h341 == io_in_csr_id ? reg_mepc : _io_out_r_csr_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_out_r_csr_T_5 = 32'h342 == io_in_csr_id ? reg_mcause : _io_out_r_csr_T_3; // @[Mux.scala 81:58]
  assign io_out_csr_br = 3'h2 == io_in_op | 3'h1 == io_in_op; // @[Mux.scala 81:58]
  assign io_out_csr_addr = 3'h2 == io_in_op ? reg_mepc : _io_out_csr_addr_T_1; // @[Mux.scala 81:58]
  assign io_out_r_csr = 32'h300 == io_in_csr_id ? reg_mstatus : _io_out_r_csr_T_5; // @[Mux.scala 81:58]
  assign io_out_difftest_mcause = reg_mcause; // @[csr.scala 125:27]
  assign io_out_difftest_mepc = reg_mepc; // @[csr.scala 126:27]
  assign io_out_difftest_mstatus = reg_mstatus; // @[csr.scala 127:27]
  assign io_out_difftest_mtvec = reg_mtvec; // @[csr.scala 128:27]
  always @(posedge clock) begin
    if (reset) begin // @[csr.scala 32:28]
      reg_mepc <= 32'h0; // @[csr.scala 32:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h341 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mepc <= _reg_mepc_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h341 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mepc <= io_in_wdata;
      end
    end else if (3'h1 == io_in_op) begin // @[Mux.scala 81:58]
      reg_mepc <= io_in_cur_pc;
    end
    if (reset) begin // @[csr.scala 33:28]
      reg_mcause <= 32'h0; // @[csr.scala 33:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h342 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mcause <= _reg_mcause_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h342 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mcause <= io_in_wdata;
      end
    end else if (3'h1 == io_in_op) begin // @[Mux.scala 81:58]
      reg_mcause <= 32'hb;
    end
    if (reset) begin // @[csr.scala 34:28]
      reg_mstatus <= 32'h0; // @[csr.scala 34:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h300 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mstatus <= _reg_mstatus_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h300 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mstatus <= io_in_wdata;
      end
    end else if (3'h2 == io_in_op) begin // @[Mux.scala 81:58]
      reg_mstatus <= {{1'd0}, _reg_mstatus_T_11};
    end else begin
      reg_mstatus <= _reg_mstatus_T_13;
    end
    if (reset) begin // @[csr.scala 35:28]
      reg_mtvec <= 32'h0; // @[csr.scala 35:28]
    end else if (3'h4 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h305 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mtvec <= _reg_mtvec_csrrs_T;
      end
    end else if (3'h3 == io_in_op) begin // @[Mux.scala 81:58]
      if (32'h305 == io_in_csr_id) begin // @[Mux.scala 81:58]
        reg_mtvec <= io_in_wdata;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mepc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mcause = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_mtvec = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ebreak_moudle(
  input   is_ebreak
);
  wire  EbreakBB_i1_is_ebreak; // @[ebreak.scala 21:29]
  EbreakBB EbreakBB_i1 ( // @[ebreak.scala 21:29]
    .is_ebreak(EbreakBB_i1_is_ebreak)
  );
  assign EbreakBB_i1_is_ebreak = is_ebreak; // @[ebreak.scala 23:30]
endmodule
module not_impl_moudle(
  input   not_impl
);
  wire  NotImplBB_i1_not_impl; // @[not_impl.scala 21:30]
  NotImplBB NotImplBB_i1 ( // @[not_impl.scala 21:30]
    .not_impl(NotImplBB_i1_not_impl)
  );
  assign NotImplBB_i1_not_impl = not_impl; // @[not_impl.scala 23:30]
endmodule
module EXU(
  input         clock,
  input         reset,
  output        from_ISU_ready,
  input         from_ISU_valid,
  input  [31:0] from_ISU_bits_imm,
  input  [31:0] from_ISU_bits_pc,
  input  [31:0] from_ISU_bits_rdata1,
  input  [31:0] from_ISU_bits_rdata2,
  input  [4:0]  from_ISU_bits_rd,
  input         from_ISU_bits_ctrl_sig_reg_wen,
  input  [2:0]  from_ISU_bits_ctrl_sig_fu_op,
  input         from_ISU_bits_ctrl_sig_mem_wen,
  input         from_ISU_bits_ctrl_sig_is_ebreak,
  input         from_ISU_bits_ctrl_sig_not_impl,
  input  [1:0]  from_ISU_bits_ctrl_sig_src1_op,
  input  [1:0]  from_ISU_bits_ctrl_sig_src2_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_alu_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_lsu_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_bru_op,
  input  [2:0]  from_ISU_bits_ctrl_sig_csr_op,
  input  [3:0]  from_ISU_bits_ctrl_sig_mdu_op,
  output        to_WBU_valid,
  output [31:0] to_WBU_bits_alu_result,
  output [31:0] to_WBU_bits_mdu_result,
  output [31:0] to_WBU_bits_lsu_rdata,
  output [31:0] to_WBU_bits_csr_rdata,
  output [31:0] to_WBU_bits_pc,
  output        to_WBU_bits_reg_wen,
  output [4:0]  to_WBU_bits_rd,
  output [2:0]  to_WBU_bits_fu_op,
  output        to_IFU_bits_bru_ctrl_br,
  output [31:0] to_IFU_bits_bru_addr,
  output        to_IFU_bits_csr_ctrl_br,
  output [31:0] to_IFU_bits_csr_addr,
  output [31:0] difftest_mcause,
  output [31:0] difftest_mepc,
  output [31:0] difftest_mstatus,
  output [31:0] difftest_mtvec,
  input         lsu_axi_master_ar_ready,
  output        lsu_axi_master_ar_valid,
  output [31:0] lsu_axi_master_ar_bits_addr,
  output        lsu_axi_master_r_ready,
  input         lsu_axi_master_r_valid,
  input  [31:0] lsu_axi_master_r_bits_data,
  input         lsu_axi_master_aw_ready,
  output        lsu_axi_master_aw_valid,
  output [31:0] lsu_axi_master_aw_bits_addr,
  input         lsu_axi_master_w_ready,
  output        lsu_axi_master_w_valid,
  output [31:0] lsu_axi_master_w_bits_data,
  output [3:0]  lsu_axi_master_w_bits_strb,
  output        lsu_axi_master_b_ready,
  input         lsu_axi_master_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] Alu_i_io_in_src1; // @[EXU.scala 22:37]
  wire [31:0] Alu_i_io_in_src2; // @[EXU.scala 22:37]
  wire [3:0] Alu_i_io_in_op; // @[EXU.scala 22:37]
  wire [31:0] Alu_i_io_out_result; // @[EXU.scala 22:37]
  wire [31:0] Mdu_i_io_in_src1; // @[EXU.scala 23:37]
  wire [31:0] Mdu_i_io_in_src2; // @[EXU.scala 23:37]
  wire [3:0] Mdu_i_io_in_op; // @[EXU.scala 23:37]
  wire [31:0] Mdu_i_io_out_result; // @[EXU.scala 23:37]
  wire [31:0] Bru_i_io_in_src1; // @[EXU.scala 24:37]
  wire [31:0] Bru_i_io_in_src2; // @[EXU.scala 24:37]
  wire [3:0] Bru_i_io_in_op; // @[EXU.scala 24:37]
  wire  Bru_i_io_out_ctrl_br; // @[EXU.scala 24:37]
  wire  Lsu_i_clock; // @[EXU.scala 25:37]
  wire  Lsu_i_reset; // @[EXU.scala 25:37]
  wire  Lsu_i_io_in_valid; // @[EXU.scala 25:37]
  wire  Lsu_i_io_in_mem_wen; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_io_in_addr; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_io_in_wdata; // @[EXU.scala 25:37]
  wire [3:0] Lsu_i_io_in_op; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_io_out_rdata; // @[EXU.scala 25:37]
  wire  Lsu_i_io_out_end; // @[EXU.scala 25:37]
  wire  Lsu_i_io_out_idle; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_ar_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_ar_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_ar_bits_addr; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_r_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_r_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_r_bits_data; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_aw_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_aw_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_aw_bits_addr; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_w_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_w_valid; // @[EXU.scala 25:37]
  wire [31:0] Lsu_i_axi_w_bits_data; // @[EXU.scala 25:37]
  wire [3:0] Lsu_i_axi_w_bits_strb; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_b_ready; // @[EXU.scala 25:37]
  wire  Lsu_i_axi_b_valid; // @[EXU.scala 25:37]
  wire  Csr_i_clock; // @[EXU.scala 26:37]
  wire  Csr_i_reset; // @[EXU.scala 26:37]
  wire [2:0] Csr_i_io_in_op; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_in_cur_pc; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_in_csr_id; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_in_wdata; // @[EXU.scala 26:37]
  wire  Csr_i_io_out_csr_br; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_csr_addr; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_r_csr; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mcause; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mepc; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mstatus; // @[EXU.scala 26:37]
  wire [31:0] Csr_i_io_out_difftest_mtvec; // @[EXU.scala 26:37]
  wire  ebreak_moudle_i_is_ebreak; // @[EXU.scala 27:37]
  wire  not_impl_moudle_i_not_impl; // @[EXU.scala 28:37]
  reg [1:0] state; // @[EXU.scala 37:24]
  wire  _state_T = from_ISU_ready & from_ISU_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_T_2 = Lsu_i_io_out_idle ? 2'h2 : 2'h1; // @[EXU.scala 45:29]
  wire [1:0] _state_T_3 = Lsu_i_io_out_end ? 2'h3 : 2'h2; // @[EXU.scala 51:25]
  wire [1:0] _GEN_1 = 2'h3 == state ? 2'h0 : state; // @[EXU.scala 38:20 54:19 37:24]
  wire [31:0] _Alu_i_io_in_src1_T_1 = 2'h2 == from_ISU_bits_ctrl_sig_src1_op ? from_ISU_bits_rdata1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _Alu_i_io_in_src2_T_1 = 2'h2 == from_ISU_bits_ctrl_sig_src2_op ? from_ISU_bits_rdata2 : 32'h0; // @[Mux.scala 81:58]
  Alu Alu_i ( // @[EXU.scala 22:37]
    .io_in_src1(Alu_i_io_in_src1),
    .io_in_src2(Alu_i_io_in_src2),
    .io_in_op(Alu_i_io_in_op),
    .io_out_result(Alu_i_io_out_result)
  );
  Mdu Mdu_i ( // @[EXU.scala 23:37]
    .io_in_src1(Mdu_i_io_in_src1),
    .io_in_src2(Mdu_i_io_in_src2),
    .io_in_op(Mdu_i_io_in_op),
    .io_out_result(Mdu_i_io_out_result)
  );
  Bru Bru_i ( // @[EXU.scala 24:37]
    .io_in_src1(Bru_i_io_in_src1),
    .io_in_src2(Bru_i_io_in_src2),
    .io_in_op(Bru_i_io_in_op),
    .io_out_ctrl_br(Bru_i_io_out_ctrl_br)
  );
  Lsu Lsu_i ( // @[EXU.scala 25:37]
    .clock(Lsu_i_clock),
    .reset(Lsu_i_reset),
    .io_in_valid(Lsu_i_io_in_valid),
    .io_in_mem_wen(Lsu_i_io_in_mem_wen),
    .io_in_addr(Lsu_i_io_in_addr),
    .io_in_wdata(Lsu_i_io_in_wdata),
    .io_in_op(Lsu_i_io_in_op),
    .io_out_rdata(Lsu_i_io_out_rdata),
    .io_out_end(Lsu_i_io_out_end),
    .io_out_idle(Lsu_i_io_out_idle),
    .axi_ar_ready(Lsu_i_axi_ar_ready),
    .axi_ar_valid(Lsu_i_axi_ar_valid),
    .axi_ar_bits_addr(Lsu_i_axi_ar_bits_addr),
    .axi_r_ready(Lsu_i_axi_r_ready),
    .axi_r_valid(Lsu_i_axi_r_valid),
    .axi_r_bits_data(Lsu_i_axi_r_bits_data),
    .axi_aw_ready(Lsu_i_axi_aw_ready),
    .axi_aw_valid(Lsu_i_axi_aw_valid),
    .axi_aw_bits_addr(Lsu_i_axi_aw_bits_addr),
    .axi_w_ready(Lsu_i_axi_w_ready),
    .axi_w_valid(Lsu_i_axi_w_valid),
    .axi_w_bits_data(Lsu_i_axi_w_bits_data),
    .axi_w_bits_strb(Lsu_i_axi_w_bits_strb),
    .axi_b_ready(Lsu_i_axi_b_ready),
    .axi_b_valid(Lsu_i_axi_b_valid)
  );
  Csr Csr_i ( // @[EXU.scala 26:37]
    .clock(Csr_i_clock),
    .reset(Csr_i_reset),
    .io_in_op(Csr_i_io_in_op),
    .io_in_cur_pc(Csr_i_io_in_cur_pc),
    .io_in_csr_id(Csr_i_io_in_csr_id),
    .io_in_wdata(Csr_i_io_in_wdata),
    .io_out_csr_br(Csr_i_io_out_csr_br),
    .io_out_csr_addr(Csr_i_io_out_csr_addr),
    .io_out_r_csr(Csr_i_io_out_r_csr),
    .io_out_difftest_mcause(Csr_i_io_out_difftest_mcause),
    .io_out_difftest_mepc(Csr_i_io_out_difftest_mepc),
    .io_out_difftest_mstatus(Csr_i_io_out_difftest_mstatus),
    .io_out_difftest_mtvec(Csr_i_io_out_difftest_mtvec)
  );
  ebreak_moudle ebreak_moudle_i ( // @[EXU.scala 27:37]
    .is_ebreak(ebreak_moudle_i_is_ebreak)
  );
  not_impl_moudle not_impl_moudle_i ( // @[EXU.scala 28:37]
    .not_impl(not_impl_moudle_i_not_impl)
  );
  assign from_ISU_ready = 2'h0 == state; // @[Mux.scala 81:61]
  assign to_WBU_valid = 2'h3 == state; // @[Mux.scala 81:61]
  assign to_WBU_bits_alu_result = Alu_i_io_out_result; // @[EXU.scala 102:28]
  assign to_WBU_bits_mdu_result = Mdu_i_io_out_result; // @[EXU.scala 103:28]
  assign to_WBU_bits_lsu_rdata = Lsu_i_io_out_rdata; // @[EXU.scala 104:28]
  assign to_WBU_bits_csr_rdata = Csr_i_io_out_r_csr; // @[EXU.scala 105:28]
  assign to_WBU_bits_pc = from_ISU_bits_pc; // @[EXU.scala 107:28]
  assign to_WBU_bits_reg_wen = from_ISU_bits_ctrl_sig_reg_wen; // @[EXU.scala 108:28]
  assign to_WBU_bits_rd = from_ISU_bits_rd; // @[EXU.scala 110:28]
  assign to_WBU_bits_fu_op = from_ISU_bits_ctrl_sig_fu_op; // @[EXU.scala 109:28]
  assign to_IFU_bits_bru_ctrl_br = Bru_i_io_out_ctrl_br; // @[EXU.scala 112:33]
  assign to_IFU_bits_bru_addr = Alu_i_io_out_result; // @[EXU.scala 113:33]
  assign to_IFU_bits_csr_ctrl_br = Csr_i_io_out_csr_br; // @[EXU.scala 114:33]
  assign to_IFU_bits_csr_addr = Csr_i_io_out_csr_addr; // @[EXU.scala 115:33]
  assign difftest_mcause = Csr_i_io_out_difftest_mcause; // @[EXU.scala 117:14]
  assign difftest_mepc = Csr_i_io_out_difftest_mepc; // @[EXU.scala 117:14]
  assign difftest_mstatus = Csr_i_io_out_difftest_mstatus; // @[EXU.scala 117:14]
  assign difftest_mtvec = Csr_i_io_out_difftest_mtvec; // @[EXU.scala 117:14]
  assign lsu_axi_master_ar_valid = Lsu_i_axi_ar_valid; // @[EXU.scala 118:20]
  assign lsu_axi_master_ar_bits_addr = Lsu_i_axi_ar_bits_addr; // @[EXU.scala 118:20]
  assign lsu_axi_master_r_ready = Lsu_i_axi_r_ready; // @[EXU.scala 118:20]
  assign lsu_axi_master_aw_valid = Lsu_i_axi_aw_valid; // @[EXU.scala 118:20]
  assign lsu_axi_master_aw_bits_addr = Lsu_i_axi_aw_bits_addr; // @[EXU.scala 118:20]
  assign lsu_axi_master_w_valid = Lsu_i_axi_w_valid; // @[EXU.scala 118:20]
  assign lsu_axi_master_w_bits_data = Lsu_i_axi_w_bits_data; // @[EXU.scala 118:20]
  assign lsu_axi_master_w_bits_strb = Lsu_i_axi_w_bits_strb; // @[EXU.scala 118:20]
  assign lsu_axi_master_b_ready = Lsu_i_axi_b_ready; // @[EXU.scala 118:20]
  assign Alu_i_io_in_src1 = 2'h1 == from_ISU_bits_ctrl_sig_src1_op ? from_ISU_bits_pc : _Alu_i_io_in_src1_T_1; // @[Mux.scala 81:58]
  assign Alu_i_io_in_src2 = 2'h3 == from_ISU_bits_ctrl_sig_src2_op ? from_ISU_bits_imm : _Alu_i_io_in_src2_T_1; // @[Mux.scala 81:58]
  assign Alu_i_io_in_op = from_ISU_bits_ctrl_sig_alu_op; // @[EXU.scala 62:20]
  assign Mdu_i_io_in_src1 = from_ISU_bits_rdata1; // @[EXU.scala 74:24]
  assign Mdu_i_io_in_src2 = from_ISU_bits_rdata2; // @[EXU.scala 75:24]
  assign Mdu_i_io_in_op = from_ISU_bits_ctrl_sig_mdu_op; // @[EXU.scala 73:24]
  assign Bru_i_io_in_src1 = from_ISU_bits_rdata1; // @[EXU.scala 87:24]
  assign Bru_i_io_in_src2 = from_ISU_bits_rdata2; // @[EXU.scala 88:24]
  assign Bru_i_io_in_op = from_ISU_bits_ctrl_sig_bru_op; // @[EXU.scala 86:24]
  assign Lsu_i_clock = clock;
  assign Lsu_i_reset = reset;
  assign Lsu_i_io_in_valid = 2'h2 == state; // @[Mux.scala 81:61]
  assign Lsu_i_io_in_mem_wen = from_ISU_bits_ctrl_sig_mem_wen; // @[EXU.scala 80:25]
  assign Lsu_i_io_in_addr = Alu_i_io_out_result; // @[EXU.scala 78:25]
  assign Lsu_i_io_in_wdata = from_ISU_bits_rdata2; // @[EXU.scala 79:25]
  assign Lsu_i_io_in_op = from_ISU_bits_ctrl_sig_lsu_op; // @[EXU.scala 81:25]
  assign Lsu_i_axi_ar_ready = lsu_axi_master_ar_ready; // @[EXU.scala 118:20]
  assign Lsu_i_axi_r_valid = lsu_axi_master_r_valid; // @[EXU.scala 118:20]
  assign Lsu_i_axi_r_bits_data = lsu_axi_master_r_bits_data; // @[EXU.scala 118:20]
  assign Lsu_i_axi_aw_ready = lsu_axi_master_aw_ready; // @[EXU.scala 118:20]
  assign Lsu_i_axi_w_ready = lsu_axi_master_w_ready; // @[EXU.scala 118:20]
  assign Lsu_i_axi_b_valid = lsu_axi_master_b_valid; // @[EXU.scala 118:20]
  assign Csr_i_clock = clock;
  assign Csr_i_reset = reset;
  assign Csr_i_io_in_op = from_ISU_bits_ctrl_sig_csr_op; // @[EXU.scala 91:25]
  assign Csr_i_io_in_cur_pc = from_ISU_bits_pc; // @[EXU.scala 92:25]
  assign Csr_i_io_in_csr_id = from_ISU_bits_imm; // @[EXU.scala 93:25]
  assign Csr_i_io_in_wdata = from_ISU_bits_rdata1; // @[EXU.scala 95:25]
  assign ebreak_moudle_i_is_ebreak = from_ISU_bits_ctrl_sig_is_ebreak; // @[EXU.scala 98:32]
  assign not_impl_moudle_i_not_impl = from_ISU_bits_ctrl_sig_not_impl; // @[EXU.scala 100:32]
  always @(posedge clock) begin
    if (reset) begin // @[EXU.scala 37:24]
      state <= 2'h0; // @[EXU.scala 37:24]
    end else if (2'h0 == state) begin // @[EXU.scala 38:20]
      if (_state_T) begin // @[EXU.scala 40:25]
        state <= 2'h1;
      end else begin
        state <= 2'h0;
      end
    end else if (2'h1 == state) begin // @[EXU.scala 38:20]
      if (from_ISU_bits_ctrl_sig_fu_op == 3'h4) begin // @[EXU.scala 44:69]
        state <= _state_T_2; // @[EXU.scala 45:23]
      end else begin
        state <= 2'h3; // @[EXU.scala 47:23]
      end
    end else if (2'h2 == state) begin // @[EXU.scala 38:20]
      state <= _state_T_3; // @[EXU.scala 51:19]
    end else begin
      state <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  output        from_EXU_ready,
  input         from_EXU_valid,
  input  [31:0] from_EXU_bits_alu_result,
  input  [31:0] from_EXU_bits_mdu_result,
  input  [31:0] from_EXU_bits_lsu_rdata,
  input  [31:0] from_EXU_bits_csr_rdata,
  input  [31:0] from_EXU_bits_pc,
  input         from_EXU_bits_reg_wen,
  input  [4:0]  from_EXU_bits_rd,
  input  [2:0]  from_EXU_bits_fu_op,
  output        to_ISU_bits_reg_wen,
  output [31:0] to_ISU_bits_wdata,
  output [4:0]  to_ISU_bits_rd,
  output        to_IFU_valid
);
  wire  _to_ISU_bits_reg_wen_T = from_EXU_ready & from_EXU_valid; // @[Decoupled.scala 51:35]
  wire [31:0] _to_ISU_bits_wdata_T_1 = from_EXU_bits_pc + 32'h4; // @[WBU.scala 25:47]
  wire [31:0] _to_ISU_bits_wdata_T_3 = 3'h1 == from_EXU_bits_fu_op ? from_EXU_bits_alu_result : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_wdata_T_5 = 3'h4 == from_EXU_bits_fu_op ? from_EXU_bits_lsu_rdata : _to_ISU_bits_wdata_T_3; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_wdata_T_7 = 3'h3 == from_EXU_bits_fu_op ? _to_ISU_bits_wdata_T_1 : _to_ISU_bits_wdata_T_5; // @[Mux.scala 81:58]
  wire [31:0] _to_ISU_bits_wdata_T_9 = 3'h5 == from_EXU_bits_fu_op ? from_EXU_bits_csr_rdata : _to_ISU_bits_wdata_T_7; // @[Mux.scala 81:58]
  assign from_EXU_ready = 1'h1; // @[WBU.scala 14:20]
  assign to_ISU_bits_reg_wen = _to_ISU_bits_reg_wen_T & from_EXU_bits_reg_wen; // @[WBU.scala 19:31]
  assign to_ISU_bits_wdata = 3'h2 == from_EXU_bits_fu_op ? from_EXU_bits_mdu_result : _to_ISU_bits_wdata_T_9; // @[Mux.scala 81:58]
  assign to_ISU_bits_rd = from_EXU_bits_rd; // @[WBU.scala 20:25]
  assign to_IFU_valid = from_EXU_valid; // @[WBU.scala 16:20]
endmodule
module IFU_cache(
  input         clock,
  input         reset,
  output        to_IDU_valid,
  output [31:0] to_IDU_bits_inst,
  output [31:0] to_IDU_bits_pc,
  input         from_EXU_bits_bru_ctrl_br,
  input  [31:0] from_EXU_bits_bru_addr,
  input         from_EXU_bits_csr_ctrl_br,
  input  [31:0] from_EXU_bits_csr_addr,
  output        from_WBU_ready,
  input         from_WBU_valid,
  input         to_cache_ready,
  output        to_cache_valid,
  output [31:0] to_cache_bits_addr,
  output        from_cache_ready,
  input         from_cache_valid,
  input  [31:0] from_cache_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_PC; // @[IFU.scala 148:26]
  wire [31:0] _next_PC_T_1 = reg_PC + 32'h4; // @[IFU.scala 156:27]
  wire  _reg_PC_T = from_WBU_ready & from_WBU_valid; // @[Decoupled.scala 51:35]
  reg [1:0] state_ifu; // @[IFU.scala 164:28]
  wire  _state_ifu_T = to_cache_ready & to_cache_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_ifu_T_1 = _state_ifu_T ? 2'h1 : 2'h0; // @[IFU.scala 166:26]
  wire  _state_ifu_T_2 = from_cache_ready & from_cache_valid; // @[Decoupled.scala 51:35]
  assign to_IDU_valid = 2'h2 == state_ifu; // @[Mux.scala 81:61]
  assign to_IDU_bits_inst = to_IDU_valid ? from_cache_bits_data : 32'h13; // @[IFU.scala 178:28]
  assign to_IDU_bits_pc = reg_PC; // @[IFU.scala 179:22]
  assign from_WBU_ready = 2'h2 == state_ifu; // @[Mux.scala 81:61]
  assign to_cache_valid = 2'h0 == state_ifu; // @[Mux.scala 81:61]
  assign to_cache_bits_addr = reg_PC; // @[IFU.scala 173:24]
  assign from_cache_ready = 2'h1 == state_ifu; // @[Mux.scala 81:61]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 148:26]
      reg_PC <= 32'h80000000; // @[IFU.scala 148:26]
    end else if (_reg_PC_T) begin // @[IFU.scala 160:18]
      if (from_EXU_bits_bru_ctrl_br) begin // @[IFU.scala 151:38]
        reg_PC <= from_EXU_bits_bru_addr; // @[IFU.scala 152:17]
      end else if (from_EXU_bits_csr_ctrl_br) begin // @[IFU.scala 153:45]
        reg_PC <= from_EXU_bits_csr_addr; // @[IFU.scala 154:17]
      end else begin
        reg_PC <= _next_PC_T_1; // @[IFU.scala 156:17]
      end
    end
    if (reset) begin // @[IFU.scala 164:28]
      state_ifu <= 2'h0; // @[IFU.scala 164:28]
    end else if (2'h2 == state_ifu) begin // @[Mux.scala 81:58]
      if (_reg_PC_T) begin // @[IFU.scala 168:28]
        state_ifu <= 2'h0;
      end else begin
        state_ifu <= 2'h2;
      end
    end else if (2'h1 == state_ifu) begin // @[Mux.scala 81:58]
      if (_state_ifu_T_2) begin // @[IFU.scala 167:28]
        state_ifu <= 2'h2;
      end else begin
        state_ifu <= 2'h1;
      end
    end else if (2'h0 == state_ifu) begin // @[Mux.scala 81:58]
      state_ifu <= _state_ifu_T_1;
    end else begin
      state_ifu <= 2'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_PC = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  state_ifu = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module I_Cache(
  input         clock,
  input         reset,
  output        from_IFU_ready,
  input         from_IFU_valid,
  input  [31:0] from_IFU_bits_addr,
  output        to_IFU_valid,
  output [31:0] to_IFU_bits_data,
  input         to_sram_ar_ready,
  output        to_sram_ar_valid,
  output [31:0] to_sram_ar_bits_addr,
  output [7:0]  to_sram_ar_bits_len,
  output        to_sram_r_ready,
  input         to_sram_r_valid,
  input  [31:0] to_sram_r_bits_data,
  input         to_sram_r_bits_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_765;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] dataArray_0_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_0_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_0_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_0_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_0_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_0_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_0_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_0_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_0_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_0_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_1_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_1_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_1_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_1_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_1_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_1_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_1_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_1_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_1_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_2_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_2_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_2_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_2_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_2_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_2_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_2_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_2_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_2_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_3_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_3_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_3_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_3_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_3_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_3_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_3_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_3_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_3_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_4_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_4_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_4_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_4_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_4_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_4_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_4_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_4_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_4_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_5_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_5_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_5_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_5_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_5_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_5_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_5_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_5_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_5_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_6_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_6_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_6_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_6_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_6_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_6_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_6_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_6_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_6_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_7_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_7_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_7_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_7_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_7_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_7_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_7_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_7_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_7_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_8_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_8_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_8_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_8_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_8_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_8_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_8_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_8_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_8_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_9_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_9_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_9_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_9_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_9_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_9_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_9_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_9_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_9_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_10_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_10_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_10_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_10_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_10_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_10_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_10_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_10_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_10_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_11_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_11_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_11_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_11_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_11_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_11_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_11_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_11_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_11_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_12_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_12_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_12_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_12_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_12_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_12_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_12_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_12_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_12_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_13_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_13_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_13_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_13_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_13_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_13_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_13_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_13_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_13_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_14_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_14_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_14_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_14_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_14_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_14_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_14_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_14_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_14_15_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_0 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_0_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_0_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_0_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_0_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_0_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_0_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_0_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_0_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_0_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_1 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_1_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_1_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_1_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_1_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_1_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_1_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_1_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_1_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_1_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_2 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_2_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_2_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_2_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_2_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_2_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_2_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_2_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_2_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_2_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_3 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_3_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_3_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_3_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_3_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_3_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_3_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_3_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_3_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_3_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_4 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_4_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_4_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_4_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_4_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_4_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_4_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_4_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_4_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_4_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_5 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_5_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_5_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_5_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_5_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_5_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_5_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_5_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_5_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_5_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_6 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_6_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_6_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_6_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_6_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_6_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_6_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_6_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_6_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_6_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_7 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_7_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_7_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_7_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_7_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_7_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_7_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_7_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_7_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_7_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_8 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_8_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_8_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_8_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_8_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_8_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_8_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_8_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_8_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_8_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_9 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_9_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_9_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_9_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_9_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_9_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_9_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_9_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_9_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_9_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_10 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_10_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_10_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_10_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_10_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_10_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_10_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_10_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_10_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_10_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_11 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_11_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_11_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_11_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_11_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_11_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_11_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_11_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_11_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_11_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_12 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_12_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_12_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_12_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_12_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_12_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_12_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_12_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_12_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_12_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_13 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_13_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_13_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_13_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_13_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_13_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_13_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_13_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_13_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_13_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_14 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_14_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_14_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_14_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_14_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_14_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_14_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_14_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_14_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_14_cachedata_MPORT_addr_pipe_0;
  reg [31:0] dataArray_15_15 [0:1]; // @[cache.scala 30:33]
  wire  dataArray_15_15_cachedata_MPORT_en; // @[cache.scala 30:33]
  wire  dataArray_15_15_cachedata_MPORT_addr; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_15_cachedata_MPORT_data; // @[cache.scala 30:33]
  wire [31:0] dataArray_15_15_MPORT_data; // @[cache.scala 30:33]
  wire  dataArray_15_15_MPORT_addr; // @[cache.scala 30:33]
  wire  dataArray_15_15_MPORT_mask; // @[cache.scala 30:33]
  wire  dataArray_15_15_MPORT_en; // @[cache.scala 30:33]
  reg  dataArray_15_15_cachedata_MPORT_en_pipe_0;
  reg  dataArray_15_15_cachedata_MPORT_addr_pipe_0;
  reg  replace_set; // @[cache.scala 21:30]
  wire [5:0] EntId = from_IFU_bits_addr[5:0] / 3'h4; // @[cache.scala 22:59]
  wire [3:0] CacheLineId = from_IFU_bits_addr[9:6]; // @[cache.scala 23:41]
  wire [21:0] tag = from_IFU_bits_addr[31:10]; // @[cache.scala 24:39]
  reg  random_num; // @[cache.scala 27:29]
  reg [21:0] tagArray_0_0; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_1; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_2; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_3; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_4; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_5; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_6; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_7; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_8; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_9; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_10; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_11; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_12; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_13; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_14; // @[cache.scala 31:29]
  reg [21:0] tagArray_0_15; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_0; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_1; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_2; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_3; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_4; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_5; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_6; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_7; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_8; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_9; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_10; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_11; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_12; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_13; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_14; // @[cache.scala 31:29]
  reg [21:0] tagArray_1_15; // @[cache.scala 31:29]
  reg  validArray_0_0; // @[cache.scala 32:29]
  reg  validArray_0_1; // @[cache.scala 32:29]
  reg  validArray_0_2; // @[cache.scala 32:29]
  reg  validArray_0_3; // @[cache.scala 32:29]
  reg  validArray_0_4; // @[cache.scala 32:29]
  reg  validArray_0_5; // @[cache.scala 32:29]
  reg  validArray_0_6; // @[cache.scala 32:29]
  reg  validArray_0_7; // @[cache.scala 32:29]
  reg  validArray_0_8; // @[cache.scala 32:29]
  reg  validArray_0_9; // @[cache.scala 32:29]
  reg  validArray_0_10; // @[cache.scala 32:29]
  reg  validArray_0_11; // @[cache.scala 32:29]
  reg  validArray_0_12; // @[cache.scala 32:29]
  reg  validArray_0_13; // @[cache.scala 32:29]
  reg  validArray_0_14; // @[cache.scala 32:29]
  reg  validArray_0_15; // @[cache.scala 32:29]
  reg  validArray_1_0; // @[cache.scala 32:29]
  reg  validArray_1_1; // @[cache.scala 32:29]
  reg  validArray_1_2; // @[cache.scala 32:29]
  reg  validArray_1_3; // @[cache.scala 32:29]
  reg  validArray_1_4; // @[cache.scala 32:29]
  reg  validArray_1_5; // @[cache.scala 32:29]
  reg  validArray_1_6; // @[cache.scala 32:29]
  reg  validArray_1_7; // @[cache.scala 32:29]
  reg  validArray_1_8; // @[cache.scala 32:29]
  reg  validArray_1_9; // @[cache.scala 32:29]
  reg  validArray_1_10; // @[cache.scala 32:29]
  reg  validArray_1_11; // @[cache.scala 32:29]
  reg  validArray_1_12; // @[cache.scala 32:29]
  reg  validArray_1_13; // @[cache.scala 32:29]
  reg  validArray_1_14; // @[cache.scala 32:29]
  reg  validArray_1_15; // @[cache.scala 32:29]
  wire [21:0] _GEN_1 = 4'h1 == CacheLineId ? tagArray_0_1 : tagArray_0_0; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_2 = 4'h2 == CacheLineId ? tagArray_0_2 : _GEN_1; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_3 = 4'h3 == CacheLineId ? tagArray_0_3 : _GEN_2; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_4 = 4'h4 == CacheLineId ? tagArray_0_4 : _GEN_3; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_5 = 4'h5 == CacheLineId ? tagArray_0_5 : _GEN_4; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_6 = 4'h6 == CacheLineId ? tagArray_0_6 : _GEN_5; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_7 = 4'h7 == CacheLineId ? tagArray_0_7 : _GEN_6; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_8 = 4'h8 == CacheLineId ? tagArray_0_8 : _GEN_7; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_9 = 4'h9 == CacheLineId ? tagArray_0_9 : _GEN_8; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_10 = 4'ha == CacheLineId ? tagArray_0_10 : _GEN_9; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_11 = 4'hb == CacheLineId ? tagArray_0_11 : _GEN_10; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_12 = 4'hc == CacheLineId ? tagArray_0_12 : _GEN_11; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_13 = 4'hd == CacheLineId ? tagArray_0_13 : _GEN_12; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_14 = 4'he == CacheLineId ? tagArray_0_14 : _GEN_13; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_15 = 4'hf == CacheLineId ? tagArray_0_15 : _GEN_14; // @[cache.scala 36:{14,14}]
  wire  _GEN_17 = 4'h1 == CacheLineId ? validArray_0_1 : validArray_0_0; // @[cache.scala 36:{44,44}]
  wire  _GEN_18 = 4'h2 == CacheLineId ? validArray_0_2 : _GEN_17; // @[cache.scala 36:{44,44}]
  wire  _GEN_19 = 4'h3 == CacheLineId ? validArray_0_3 : _GEN_18; // @[cache.scala 36:{44,44}]
  wire  _GEN_20 = 4'h4 == CacheLineId ? validArray_0_4 : _GEN_19; // @[cache.scala 36:{44,44}]
  wire  _GEN_21 = 4'h5 == CacheLineId ? validArray_0_5 : _GEN_20; // @[cache.scala 36:{44,44}]
  wire  _GEN_22 = 4'h6 == CacheLineId ? validArray_0_6 : _GEN_21; // @[cache.scala 36:{44,44}]
  wire  _GEN_23 = 4'h7 == CacheLineId ? validArray_0_7 : _GEN_22; // @[cache.scala 36:{44,44}]
  wire  _GEN_24 = 4'h8 == CacheLineId ? validArray_0_8 : _GEN_23; // @[cache.scala 36:{44,44}]
  wire  _GEN_25 = 4'h9 == CacheLineId ? validArray_0_9 : _GEN_24; // @[cache.scala 36:{44,44}]
  wire  _GEN_26 = 4'ha == CacheLineId ? validArray_0_10 : _GEN_25; // @[cache.scala 36:{44,44}]
  wire  _GEN_27 = 4'hb == CacheLineId ? validArray_0_11 : _GEN_26; // @[cache.scala 36:{44,44}]
  wire  _GEN_28 = 4'hc == CacheLineId ? validArray_0_12 : _GEN_27; // @[cache.scala 36:{44,44}]
  wire  _GEN_29 = 4'hd == CacheLineId ? validArray_0_13 : _GEN_28; // @[cache.scala 36:{44,44}]
  wire  _GEN_30 = 4'he == CacheLineId ? validArray_0_14 : _GEN_29; // @[cache.scala 36:{44,44}]
  wire  _GEN_31 = 4'hf == CacheLineId ? validArray_0_15 : _GEN_30; // @[cache.scala 36:{44,44}]
  wire  hitArray_0 = tag == _GEN_15 & _GEN_31; // @[cache.scala 36:44]
  wire [21:0] _GEN_33 = 4'h1 == CacheLineId ? tagArray_1_1 : tagArray_1_0; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_34 = 4'h2 == CacheLineId ? tagArray_1_2 : _GEN_33; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_35 = 4'h3 == CacheLineId ? tagArray_1_3 : _GEN_34; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_36 = 4'h4 == CacheLineId ? tagArray_1_4 : _GEN_35; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_37 = 4'h5 == CacheLineId ? tagArray_1_5 : _GEN_36; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_38 = 4'h6 == CacheLineId ? tagArray_1_6 : _GEN_37; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_39 = 4'h7 == CacheLineId ? tagArray_1_7 : _GEN_38; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_40 = 4'h8 == CacheLineId ? tagArray_1_8 : _GEN_39; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_41 = 4'h9 == CacheLineId ? tagArray_1_9 : _GEN_40; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_42 = 4'ha == CacheLineId ? tagArray_1_10 : _GEN_41; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_43 = 4'hb == CacheLineId ? tagArray_1_11 : _GEN_42; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_44 = 4'hc == CacheLineId ? tagArray_1_12 : _GEN_43; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_45 = 4'hd == CacheLineId ? tagArray_1_13 : _GEN_44; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_46 = 4'he == CacheLineId ? tagArray_1_14 : _GEN_45; // @[cache.scala 36:{14,14}]
  wire [21:0] _GEN_47 = 4'hf == CacheLineId ? tagArray_1_15 : _GEN_46; // @[cache.scala 36:{14,14}]
  wire  _GEN_49 = 4'h1 == CacheLineId ? validArray_1_1 : validArray_1_0; // @[cache.scala 36:{44,44}]
  wire  _GEN_50 = 4'h2 == CacheLineId ? validArray_1_2 : _GEN_49; // @[cache.scala 36:{44,44}]
  wire  _GEN_51 = 4'h3 == CacheLineId ? validArray_1_3 : _GEN_50; // @[cache.scala 36:{44,44}]
  wire  _GEN_52 = 4'h4 == CacheLineId ? validArray_1_4 : _GEN_51; // @[cache.scala 36:{44,44}]
  wire  _GEN_53 = 4'h5 == CacheLineId ? validArray_1_5 : _GEN_52; // @[cache.scala 36:{44,44}]
  wire  _GEN_54 = 4'h6 == CacheLineId ? validArray_1_6 : _GEN_53; // @[cache.scala 36:{44,44}]
  wire  _GEN_55 = 4'h7 == CacheLineId ? validArray_1_7 : _GEN_54; // @[cache.scala 36:{44,44}]
  wire  _GEN_56 = 4'h8 == CacheLineId ? validArray_1_8 : _GEN_55; // @[cache.scala 36:{44,44}]
  wire  _GEN_57 = 4'h9 == CacheLineId ? validArray_1_9 : _GEN_56; // @[cache.scala 36:{44,44}]
  wire  _GEN_58 = 4'ha == CacheLineId ? validArray_1_10 : _GEN_57; // @[cache.scala 36:{44,44}]
  wire  _GEN_59 = 4'hb == CacheLineId ? validArray_1_11 : _GEN_58; // @[cache.scala 36:{44,44}]
  wire  _GEN_60 = 4'hc == CacheLineId ? validArray_1_12 : _GEN_59; // @[cache.scala 36:{44,44}]
  wire  _GEN_61 = 4'hd == CacheLineId ? validArray_1_13 : _GEN_60; // @[cache.scala 36:{44,44}]
  wire  _GEN_62 = 4'he == CacheLineId ? validArray_1_14 : _GEN_61; // @[cache.scala 36:{44,44}]
  wire  _GEN_63 = 4'hf == CacheLineId ? validArray_1_15 : _GEN_62; // @[cache.scala 36:{44,44}]
  wire  hitArray_1 = tag == _GEN_47 & _GEN_63; // @[cache.scala 36:44]
  wire  hit = hitArray_0 | hitArray_1; // @[cache.scala 38:33]
  reg [3:0] off; // @[cache.scala 45:24]
  reg [2:0] state_cache; // @[cache.scala 48:30]
  wire  _T_1 = from_IFU_ready & from_IFU_valid; // @[Decoupled.scala 51:35]
  wire  _T_3 = 3'h2 == state_cache; // @[cache.scala 49:26]
  wire  _state_cache_T_1 = to_sram_ar_ready & to_sram_ar_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_cache_T_2 = _state_cache_T_1 ? 3'h3 : 3'h2; // @[cache.scala 62:31]
  wire [2:0] _state_cache_T_3 = to_sram_r_bits_last ? 3'h4 : 3'h3; // @[cache.scala 68:31]
  wire  _off_T = to_sram_r_ready & to_sram_r_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _off_T_2 = off + 4'h1; // @[cache.scala 69:51]
  wire [3:0] _off_T_3 = _off_T ? _off_T_2 : off; // @[cache.scala 69:31]
  wire [2:0] _GEN_65 = 3'h4 == state_cache ? 3'h1 : state_cache; // @[cache.scala 49:26 74:25 48:30]
  wire [2:0] _GEN_66 = 3'h3 == state_cache ? _state_cache_T_3 : _GEN_65; // @[cache.scala 49:26 68:25]
  wire [3:0] _GEN_67 = 3'h3 == state_cache ? _off_T_3 : off; // @[cache.scala 45:24 49:26 69:25]
  wire  _T_6 = state_cache == 3'h3; // @[cache.scala 80:24]
  wire  _GEN_1552 = 4'h0 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1553 = 4'h0 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1555 = 4'h1 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1557 = 4'h2 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1559 = 4'h3 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1561 = 4'h4 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1563 = 4'h5 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1565 = 4'h6 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1567 = 4'h7 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1569 = 4'h8 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1571 = 4'h9 == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1573 = 4'ha == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1575 = 4'hb == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1577 = 4'hc == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1579 = 4'hd == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1581 = 4'he == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1583 = 4'hf == off; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1584 = 4'h1 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1616 = 4'h2 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1648 = 4'h3 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1680 = 4'h4 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1712 = 4'h5 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1744 = 4'h6 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1776 = 4'h7 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1808 = 4'h8 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1840 = 4'h9 == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1872 = 4'ha == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1904 = 4'hb == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1936 = 4'hc == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_1968 = 4'hd == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_2000 = 4'he == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_2032 = 4'hf == CacheLineId; // @[cache.scala 81:{18,50,50}]
  wire  _GEN_2064 = ~replace_set; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_589 = ~replace_set & _GEN_1552 | validArray_0_0; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_590 = ~replace_set & _GEN_1584 | validArray_0_1; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_591 = ~replace_set & _GEN_1616 | validArray_0_2; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_592 = ~replace_set & _GEN_1648 | validArray_0_3; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_593 = ~replace_set & _GEN_1680 | validArray_0_4; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_594 = ~replace_set & _GEN_1712 | validArray_0_5; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_595 = ~replace_set & _GEN_1744 | validArray_0_6; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_596 = ~replace_set & _GEN_1776 | validArray_0_7; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_597 = ~replace_set & _GEN_1808 | validArray_0_8; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_598 = ~replace_set & _GEN_1840 | validArray_0_9; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_599 = ~replace_set & _GEN_1872 | validArray_0_10; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_600 = ~replace_set & _GEN_1904 | validArray_0_11; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_601 = ~replace_set & _GEN_1936 | validArray_0_12; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_602 = ~replace_set & _GEN_1968 | validArray_0_13; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_603 = ~replace_set & _GEN_2000 | validArray_0_14; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_604 = ~replace_set & _GEN_2032 | validArray_0_15; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_605 = replace_set & _GEN_1552 | validArray_1_0; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_606 = replace_set & _GEN_1584 | validArray_1_1; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_607 = replace_set & _GEN_1616 | validArray_1_2; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_608 = replace_set & _GEN_1648 | validArray_1_3; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_609 = replace_set & _GEN_1680 | validArray_1_4; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_610 = replace_set & _GEN_1712 | validArray_1_5; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_611 = replace_set & _GEN_1744 | validArray_1_6; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_612 = replace_set & _GEN_1776 | validArray_1_7; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_613 = replace_set & _GEN_1808 | validArray_1_8; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_614 = replace_set & _GEN_1840 | validArray_1_9; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_615 = replace_set & _GEN_1872 | validArray_1_10; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_616 = replace_set & _GEN_1904 | validArray_1_11; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_617 = replace_set & _GEN_1936 | validArray_1_12; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_618 = replace_set & _GEN_1968 | validArray_1_13; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_619 = replace_set & _GEN_2000 | validArray_1_14; // @[cache.scala 32:29 83:{50,50}]
  wire  _GEN_620 = replace_set & _GEN_2032 | validArray_1_15; // @[cache.scala 32:29 83:{50,50}]
  wire [31:0] _to_sram_ar_bits_addr_T = {{6'd0}, from_IFU_bits_addr[31:6]}; // @[cache.scala 91:91]
  wire [37:0] _GEN_2193 = {_to_sram_ar_bits_addr_T, 6'h0}; // @[cache.scala 91:104]
  wire [38:0] _to_sram_ar_bits_addr_T_1 = {{1'd0}, _GEN_2193}; // @[cache.scala 91:104]
  wire [38:0] _to_sram_ar_bits_addr_T_3 = _T_3 ? _to_sram_ar_bits_addr_T_1 : 39'h0; // @[Mux.scala 81:58]
  wire [3:0] _to_sram_ar_bits_len_T_1 = _T_3 ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [31:0] _GEN_1296 = dataArray_0_0_cachedata_MPORT_data; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1297 = _GEN_1552 & 4'h1 == EntId[3:0] ? dataArray_0_1_cachedata_MPORT_data : _GEN_1296; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1298 = _GEN_1552 & 4'h2 == EntId[3:0] ? dataArray_0_2_cachedata_MPORT_data : _GEN_1297; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1299 = _GEN_1552 & 4'h3 == EntId[3:0] ? dataArray_0_3_cachedata_MPORT_data : _GEN_1298; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1300 = _GEN_1552 & 4'h4 == EntId[3:0] ? dataArray_0_4_cachedata_MPORT_data : _GEN_1299; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1301 = _GEN_1552 & 4'h5 == EntId[3:0] ? dataArray_0_5_cachedata_MPORT_data : _GEN_1300; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1302 = _GEN_1552 & 4'h6 == EntId[3:0] ? dataArray_0_6_cachedata_MPORT_data : _GEN_1301; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1303 = _GEN_1552 & 4'h7 == EntId[3:0] ? dataArray_0_7_cachedata_MPORT_data : _GEN_1302; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1304 = _GEN_1552 & 4'h8 == EntId[3:0] ? dataArray_0_8_cachedata_MPORT_data : _GEN_1303; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1305 = _GEN_1552 & 4'h9 == EntId[3:0] ? dataArray_0_9_cachedata_MPORT_data : _GEN_1304; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1306 = _GEN_1552 & 4'ha == EntId[3:0] ? dataArray_0_10_cachedata_MPORT_data : _GEN_1305; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1307 = _GEN_1552 & 4'hb == EntId[3:0] ? dataArray_0_11_cachedata_MPORT_data : _GEN_1306; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1308 = _GEN_1552 & 4'hc == EntId[3:0] ? dataArray_0_12_cachedata_MPORT_data : _GEN_1307; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1309 = _GEN_1552 & 4'hd == EntId[3:0] ? dataArray_0_13_cachedata_MPORT_data : _GEN_1308; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1310 = _GEN_1552 & 4'he == EntId[3:0] ? dataArray_0_14_cachedata_MPORT_data : _GEN_1309; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1311 = _GEN_1552 & 4'hf == EntId[3:0] ? dataArray_0_15_cachedata_MPORT_data : _GEN_1310; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1312 = _GEN_1584 & 4'h0 == EntId[3:0] ? dataArray_1_0_cachedata_MPORT_data : _GEN_1311; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1313 = _GEN_1584 & 4'h1 == EntId[3:0] ? dataArray_1_1_cachedata_MPORT_data : _GEN_1312; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1314 = _GEN_1584 & 4'h2 == EntId[3:0] ? dataArray_1_2_cachedata_MPORT_data : _GEN_1313; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1315 = _GEN_1584 & 4'h3 == EntId[3:0] ? dataArray_1_3_cachedata_MPORT_data : _GEN_1314; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1316 = _GEN_1584 & 4'h4 == EntId[3:0] ? dataArray_1_4_cachedata_MPORT_data : _GEN_1315; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1317 = _GEN_1584 & 4'h5 == EntId[3:0] ? dataArray_1_5_cachedata_MPORT_data : _GEN_1316; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1318 = _GEN_1584 & 4'h6 == EntId[3:0] ? dataArray_1_6_cachedata_MPORT_data : _GEN_1317; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1319 = _GEN_1584 & 4'h7 == EntId[3:0] ? dataArray_1_7_cachedata_MPORT_data : _GEN_1318; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1320 = _GEN_1584 & 4'h8 == EntId[3:0] ? dataArray_1_8_cachedata_MPORT_data : _GEN_1319; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1321 = _GEN_1584 & 4'h9 == EntId[3:0] ? dataArray_1_9_cachedata_MPORT_data : _GEN_1320; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1322 = _GEN_1584 & 4'ha == EntId[3:0] ? dataArray_1_10_cachedata_MPORT_data : _GEN_1321; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1323 = _GEN_1584 & 4'hb == EntId[3:0] ? dataArray_1_11_cachedata_MPORT_data : _GEN_1322; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1324 = _GEN_1584 & 4'hc == EntId[3:0] ? dataArray_1_12_cachedata_MPORT_data : _GEN_1323; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1325 = _GEN_1584 & 4'hd == EntId[3:0] ? dataArray_1_13_cachedata_MPORT_data : _GEN_1324; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1326 = _GEN_1584 & 4'he == EntId[3:0] ? dataArray_1_14_cachedata_MPORT_data : _GEN_1325; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1327 = _GEN_1584 & 4'hf == EntId[3:0] ? dataArray_1_15_cachedata_MPORT_data : _GEN_1326; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1328 = _GEN_1616 & 4'h0 == EntId[3:0] ? dataArray_2_0_cachedata_MPORT_data : _GEN_1327; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1329 = _GEN_1616 & 4'h1 == EntId[3:0] ? dataArray_2_1_cachedata_MPORT_data : _GEN_1328; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1330 = _GEN_1616 & 4'h2 == EntId[3:0] ? dataArray_2_2_cachedata_MPORT_data : _GEN_1329; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1331 = _GEN_1616 & 4'h3 == EntId[3:0] ? dataArray_2_3_cachedata_MPORT_data : _GEN_1330; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1332 = _GEN_1616 & 4'h4 == EntId[3:0] ? dataArray_2_4_cachedata_MPORT_data : _GEN_1331; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1333 = _GEN_1616 & 4'h5 == EntId[3:0] ? dataArray_2_5_cachedata_MPORT_data : _GEN_1332; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1334 = _GEN_1616 & 4'h6 == EntId[3:0] ? dataArray_2_6_cachedata_MPORT_data : _GEN_1333; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1335 = _GEN_1616 & 4'h7 == EntId[3:0] ? dataArray_2_7_cachedata_MPORT_data : _GEN_1334; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1336 = _GEN_1616 & 4'h8 == EntId[3:0] ? dataArray_2_8_cachedata_MPORT_data : _GEN_1335; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1337 = _GEN_1616 & 4'h9 == EntId[3:0] ? dataArray_2_9_cachedata_MPORT_data : _GEN_1336; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1338 = _GEN_1616 & 4'ha == EntId[3:0] ? dataArray_2_10_cachedata_MPORT_data : _GEN_1337; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1339 = _GEN_1616 & 4'hb == EntId[3:0] ? dataArray_2_11_cachedata_MPORT_data : _GEN_1338; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1340 = _GEN_1616 & 4'hc == EntId[3:0] ? dataArray_2_12_cachedata_MPORT_data : _GEN_1339; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1341 = _GEN_1616 & 4'hd == EntId[3:0] ? dataArray_2_13_cachedata_MPORT_data : _GEN_1340; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1342 = _GEN_1616 & 4'he == EntId[3:0] ? dataArray_2_14_cachedata_MPORT_data : _GEN_1341; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1343 = _GEN_1616 & 4'hf == EntId[3:0] ? dataArray_2_15_cachedata_MPORT_data : _GEN_1342; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1344 = _GEN_1648 & 4'h0 == EntId[3:0] ? dataArray_3_0_cachedata_MPORT_data : _GEN_1343; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1345 = _GEN_1648 & 4'h1 == EntId[3:0] ? dataArray_3_1_cachedata_MPORT_data : _GEN_1344; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1346 = _GEN_1648 & 4'h2 == EntId[3:0] ? dataArray_3_2_cachedata_MPORT_data : _GEN_1345; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1347 = _GEN_1648 & 4'h3 == EntId[3:0] ? dataArray_3_3_cachedata_MPORT_data : _GEN_1346; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1348 = _GEN_1648 & 4'h4 == EntId[3:0] ? dataArray_3_4_cachedata_MPORT_data : _GEN_1347; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1349 = _GEN_1648 & 4'h5 == EntId[3:0] ? dataArray_3_5_cachedata_MPORT_data : _GEN_1348; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1350 = _GEN_1648 & 4'h6 == EntId[3:0] ? dataArray_3_6_cachedata_MPORT_data : _GEN_1349; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1351 = _GEN_1648 & 4'h7 == EntId[3:0] ? dataArray_3_7_cachedata_MPORT_data : _GEN_1350; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1352 = _GEN_1648 & 4'h8 == EntId[3:0] ? dataArray_3_8_cachedata_MPORT_data : _GEN_1351; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1353 = _GEN_1648 & 4'h9 == EntId[3:0] ? dataArray_3_9_cachedata_MPORT_data : _GEN_1352; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1354 = _GEN_1648 & 4'ha == EntId[3:0] ? dataArray_3_10_cachedata_MPORT_data : _GEN_1353; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1355 = _GEN_1648 & 4'hb == EntId[3:0] ? dataArray_3_11_cachedata_MPORT_data : _GEN_1354; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1356 = _GEN_1648 & 4'hc == EntId[3:0] ? dataArray_3_12_cachedata_MPORT_data : _GEN_1355; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1357 = _GEN_1648 & 4'hd == EntId[3:0] ? dataArray_3_13_cachedata_MPORT_data : _GEN_1356; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1358 = _GEN_1648 & 4'he == EntId[3:0] ? dataArray_3_14_cachedata_MPORT_data : _GEN_1357; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1359 = _GEN_1648 & 4'hf == EntId[3:0] ? dataArray_3_15_cachedata_MPORT_data : _GEN_1358; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1360 = _GEN_1680 & 4'h0 == EntId[3:0] ? dataArray_4_0_cachedata_MPORT_data : _GEN_1359; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1361 = _GEN_1680 & 4'h1 == EntId[3:0] ? dataArray_4_1_cachedata_MPORT_data : _GEN_1360; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1362 = _GEN_1680 & 4'h2 == EntId[3:0] ? dataArray_4_2_cachedata_MPORT_data : _GEN_1361; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1363 = _GEN_1680 & 4'h3 == EntId[3:0] ? dataArray_4_3_cachedata_MPORT_data : _GEN_1362; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1364 = _GEN_1680 & 4'h4 == EntId[3:0] ? dataArray_4_4_cachedata_MPORT_data : _GEN_1363; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1365 = _GEN_1680 & 4'h5 == EntId[3:0] ? dataArray_4_5_cachedata_MPORT_data : _GEN_1364; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1366 = _GEN_1680 & 4'h6 == EntId[3:0] ? dataArray_4_6_cachedata_MPORT_data : _GEN_1365; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1367 = _GEN_1680 & 4'h7 == EntId[3:0] ? dataArray_4_7_cachedata_MPORT_data : _GEN_1366; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1368 = _GEN_1680 & 4'h8 == EntId[3:0] ? dataArray_4_8_cachedata_MPORT_data : _GEN_1367; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1369 = _GEN_1680 & 4'h9 == EntId[3:0] ? dataArray_4_9_cachedata_MPORT_data : _GEN_1368; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1370 = _GEN_1680 & 4'ha == EntId[3:0] ? dataArray_4_10_cachedata_MPORT_data : _GEN_1369; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1371 = _GEN_1680 & 4'hb == EntId[3:0] ? dataArray_4_11_cachedata_MPORT_data : _GEN_1370; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1372 = _GEN_1680 & 4'hc == EntId[3:0] ? dataArray_4_12_cachedata_MPORT_data : _GEN_1371; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1373 = _GEN_1680 & 4'hd == EntId[3:0] ? dataArray_4_13_cachedata_MPORT_data : _GEN_1372; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1374 = _GEN_1680 & 4'he == EntId[3:0] ? dataArray_4_14_cachedata_MPORT_data : _GEN_1373; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1375 = _GEN_1680 & 4'hf == EntId[3:0] ? dataArray_4_15_cachedata_MPORT_data : _GEN_1374; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1376 = _GEN_1712 & 4'h0 == EntId[3:0] ? dataArray_5_0_cachedata_MPORT_data : _GEN_1375; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1377 = _GEN_1712 & 4'h1 == EntId[3:0] ? dataArray_5_1_cachedata_MPORT_data : _GEN_1376; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1378 = _GEN_1712 & 4'h2 == EntId[3:0] ? dataArray_5_2_cachedata_MPORT_data : _GEN_1377; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1379 = _GEN_1712 & 4'h3 == EntId[3:0] ? dataArray_5_3_cachedata_MPORT_data : _GEN_1378; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1380 = _GEN_1712 & 4'h4 == EntId[3:0] ? dataArray_5_4_cachedata_MPORT_data : _GEN_1379; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1381 = _GEN_1712 & 4'h5 == EntId[3:0] ? dataArray_5_5_cachedata_MPORT_data : _GEN_1380; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1382 = _GEN_1712 & 4'h6 == EntId[3:0] ? dataArray_5_6_cachedata_MPORT_data : _GEN_1381; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1383 = _GEN_1712 & 4'h7 == EntId[3:0] ? dataArray_5_7_cachedata_MPORT_data : _GEN_1382; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1384 = _GEN_1712 & 4'h8 == EntId[3:0] ? dataArray_5_8_cachedata_MPORT_data : _GEN_1383; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1385 = _GEN_1712 & 4'h9 == EntId[3:0] ? dataArray_5_9_cachedata_MPORT_data : _GEN_1384; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1386 = _GEN_1712 & 4'ha == EntId[3:0] ? dataArray_5_10_cachedata_MPORT_data : _GEN_1385; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1387 = _GEN_1712 & 4'hb == EntId[3:0] ? dataArray_5_11_cachedata_MPORT_data : _GEN_1386; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1388 = _GEN_1712 & 4'hc == EntId[3:0] ? dataArray_5_12_cachedata_MPORT_data : _GEN_1387; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1389 = _GEN_1712 & 4'hd == EntId[3:0] ? dataArray_5_13_cachedata_MPORT_data : _GEN_1388; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1390 = _GEN_1712 & 4'he == EntId[3:0] ? dataArray_5_14_cachedata_MPORT_data : _GEN_1389; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1391 = _GEN_1712 & 4'hf == EntId[3:0] ? dataArray_5_15_cachedata_MPORT_data : _GEN_1390; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1392 = _GEN_1744 & 4'h0 == EntId[3:0] ? dataArray_6_0_cachedata_MPORT_data : _GEN_1391; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1393 = _GEN_1744 & 4'h1 == EntId[3:0] ? dataArray_6_1_cachedata_MPORT_data : _GEN_1392; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1394 = _GEN_1744 & 4'h2 == EntId[3:0] ? dataArray_6_2_cachedata_MPORT_data : _GEN_1393; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1395 = _GEN_1744 & 4'h3 == EntId[3:0] ? dataArray_6_3_cachedata_MPORT_data : _GEN_1394; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1396 = _GEN_1744 & 4'h4 == EntId[3:0] ? dataArray_6_4_cachedata_MPORT_data : _GEN_1395; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1397 = _GEN_1744 & 4'h5 == EntId[3:0] ? dataArray_6_5_cachedata_MPORT_data : _GEN_1396; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1398 = _GEN_1744 & 4'h6 == EntId[3:0] ? dataArray_6_6_cachedata_MPORT_data : _GEN_1397; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1399 = _GEN_1744 & 4'h7 == EntId[3:0] ? dataArray_6_7_cachedata_MPORT_data : _GEN_1398; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1400 = _GEN_1744 & 4'h8 == EntId[3:0] ? dataArray_6_8_cachedata_MPORT_data : _GEN_1399; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1401 = _GEN_1744 & 4'h9 == EntId[3:0] ? dataArray_6_9_cachedata_MPORT_data : _GEN_1400; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1402 = _GEN_1744 & 4'ha == EntId[3:0] ? dataArray_6_10_cachedata_MPORT_data : _GEN_1401; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1403 = _GEN_1744 & 4'hb == EntId[3:0] ? dataArray_6_11_cachedata_MPORT_data : _GEN_1402; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1404 = _GEN_1744 & 4'hc == EntId[3:0] ? dataArray_6_12_cachedata_MPORT_data : _GEN_1403; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1405 = _GEN_1744 & 4'hd == EntId[3:0] ? dataArray_6_13_cachedata_MPORT_data : _GEN_1404; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1406 = _GEN_1744 & 4'he == EntId[3:0] ? dataArray_6_14_cachedata_MPORT_data : _GEN_1405; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1407 = _GEN_1744 & 4'hf == EntId[3:0] ? dataArray_6_15_cachedata_MPORT_data : _GEN_1406; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1408 = _GEN_1776 & 4'h0 == EntId[3:0] ? dataArray_7_0_cachedata_MPORT_data : _GEN_1407; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1409 = _GEN_1776 & 4'h1 == EntId[3:0] ? dataArray_7_1_cachedata_MPORT_data : _GEN_1408; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1410 = _GEN_1776 & 4'h2 == EntId[3:0] ? dataArray_7_2_cachedata_MPORT_data : _GEN_1409; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1411 = _GEN_1776 & 4'h3 == EntId[3:0] ? dataArray_7_3_cachedata_MPORT_data : _GEN_1410; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1412 = _GEN_1776 & 4'h4 == EntId[3:0] ? dataArray_7_4_cachedata_MPORT_data : _GEN_1411; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1413 = _GEN_1776 & 4'h5 == EntId[3:0] ? dataArray_7_5_cachedata_MPORT_data : _GEN_1412; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1414 = _GEN_1776 & 4'h6 == EntId[3:0] ? dataArray_7_6_cachedata_MPORT_data : _GEN_1413; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1415 = _GEN_1776 & 4'h7 == EntId[3:0] ? dataArray_7_7_cachedata_MPORT_data : _GEN_1414; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1416 = _GEN_1776 & 4'h8 == EntId[3:0] ? dataArray_7_8_cachedata_MPORT_data : _GEN_1415; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1417 = _GEN_1776 & 4'h9 == EntId[3:0] ? dataArray_7_9_cachedata_MPORT_data : _GEN_1416; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1418 = _GEN_1776 & 4'ha == EntId[3:0] ? dataArray_7_10_cachedata_MPORT_data : _GEN_1417; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1419 = _GEN_1776 & 4'hb == EntId[3:0] ? dataArray_7_11_cachedata_MPORT_data : _GEN_1418; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1420 = _GEN_1776 & 4'hc == EntId[3:0] ? dataArray_7_12_cachedata_MPORT_data : _GEN_1419; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1421 = _GEN_1776 & 4'hd == EntId[3:0] ? dataArray_7_13_cachedata_MPORT_data : _GEN_1420; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1422 = _GEN_1776 & 4'he == EntId[3:0] ? dataArray_7_14_cachedata_MPORT_data : _GEN_1421; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1423 = _GEN_1776 & 4'hf == EntId[3:0] ? dataArray_7_15_cachedata_MPORT_data : _GEN_1422; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1424 = _GEN_1808 & 4'h0 == EntId[3:0] ? dataArray_8_0_cachedata_MPORT_data : _GEN_1423; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1425 = _GEN_1808 & 4'h1 == EntId[3:0] ? dataArray_8_1_cachedata_MPORT_data : _GEN_1424; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1426 = _GEN_1808 & 4'h2 == EntId[3:0] ? dataArray_8_2_cachedata_MPORT_data : _GEN_1425; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1427 = _GEN_1808 & 4'h3 == EntId[3:0] ? dataArray_8_3_cachedata_MPORT_data : _GEN_1426; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1428 = _GEN_1808 & 4'h4 == EntId[3:0] ? dataArray_8_4_cachedata_MPORT_data : _GEN_1427; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1429 = _GEN_1808 & 4'h5 == EntId[3:0] ? dataArray_8_5_cachedata_MPORT_data : _GEN_1428; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1430 = _GEN_1808 & 4'h6 == EntId[3:0] ? dataArray_8_6_cachedata_MPORT_data : _GEN_1429; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1431 = _GEN_1808 & 4'h7 == EntId[3:0] ? dataArray_8_7_cachedata_MPORT_data : _GEN_1430; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1432 = _GEN_1808 & 4'h8 == EntId[3:0] ? dataArray_8_8_cachedata_MPORT_data : _GEN_1431; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1433 = _GEN_1808 & 4'h9 == EntId[3:0] ? dataArray_8_9_cachedata_MPORT_data : _GEN_1432; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1434 = _GEN_1808 & 4'ha == EntId[3:0] ? dataArray_8_10_cachedata_MPORT_data : _GEN_1433; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1435 = _GEN_1808 & 4'hb == EntId[3:0] ? dataArray_8_11_cachedata_MPORT_data : _GEN_1434; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1436 = _GEN_1808 & 4'hc == EntId[3:0] ? dataArray_8_12_cachedata_MPORT_data : _GEN_1435; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1437 = _GEN_1808 & 4'hd == EntId[3:0] ? dataArray_8_13_cachedata_MPORT_data : _GEN_1436; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1438 = _GEN_1808 & 4'he == EntId[3:0] ? dataArray_8_14_cachedata_MPORT_data : _GEN_1437; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1439 = _GEN_1808 & 4'hf == EntId[3:0] ? dataArray_8_15_cachedata_MPORT_data : _GEN_1438; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1440 = _GEN_1840 & 4'h0 == EntId[3:0] ? dataArray_9_0_cachedata_MPORT_data : _GEN_1439; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1441 = _GEN_1840 & 4'h1 == EntId[3:0] ? dataArray_9_1_cachedata_MPORT_data : _GEN_1440; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1442 = _GEN_1840 & 4'h2 == EntId[3:0] ? dataArray_9_2_cachedata_MPORT_data : _GEN_1441; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1443 = _GEN_1840 & 4'h3 == EntId[3:0] ? dataArray_9_3_cachedata_MPORT_data : _GEN_1442; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1444 = _GEN_1840 & 4'h4 == EntId[3:0] ? dataArray_9_4_cachedata_MPORT_data : _GEN_1443; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1445 = _GEN_1840 & 4'h5 == EntId[3:0] ? dataArray_9_5_cachedata_MPORT_data : _GEN_1444; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1446 = _GEN_1840 & 4'h6 == EntId[3:0] ? dataArray_9_6_cachedata_MPORT_data : _GEN_1445; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1447 = _GEN_1840 & 4'h7 == EntId[3:0] ? dataArray_9_7_cachedata_MPORT_data : _GEN_1446; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1448 = _GEN_1840 & 4'h8 == EntId[3:0] ? dataArray_9_8_cachedata_MPORT_data : _GEN_1447; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1449 = _GEN_1840 & 4'h9 == EntId[3:0] ? dataArray_9_9_cachedata_MPORT_data : _GEN_1448; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1450 = _GEN_1840 & 4'ha == EntId[3:0] ? dataArray_9_10_cachedata_MPORT_data : _GEN_1449; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1451 = _GEN_1840 & 4'hb == EntId[3:0] ? dataArray_9_11_cachedata_MPORT_data : _GEN_1450; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1452 = _GEN_1840 & 4'hc == EntId[3:0] ? dataArray_9_12_cachedata_MPORT_data : _GEN_1451; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1453 = _GEN_1840 & 4'hd == EntId[3:0] ? dataArray_9_13_cachedata_MPORT_data : _GEN_1452; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1454 = _GEN_1840 & 4'he == EntId[3:0] ? dataArray_9_14_cachedata_MPORT_data : _GEN_1453; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1455 = _GEN_1840 & 4'hf == EntId[3:0] ? dataArray_9_15_cachedata_MPORT_data : _GEN_1454; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1456 = _GEN_1872 & 4'h0 == EntId[3:0] ? dataArray_10_0_cachedata_MPORT_data : _GEN_1455; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1457 = _GEN_1872 & 4'h1 == EntId[3:0] ? dataArray_10_1_cachedata_MPORT_data : _GEN_1456; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1458 = _GEN_1872 & 4'h2 == EntId[3:0] ? dataArray_10_2_cachedata_MPORT_data : _GEN_1457; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1459 = _GEN_1872 & 4'h3 == EntId[3:0] ? dataArray_10_3_cachedata_MPORT_data : _GEN_1458; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1460 = _GEN_1872 & 4'h4 == EntId[3:0] ? dataArray_10_4_cachedata_MPORT_data : _GEN_1459; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1461 = _GEN_1872 & 4'h5 == EntId[3:0] ? dataArray_10_5_cachedata_MPORT_data : _GEN_1460; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1462 = _GEN_1872 & 4'h6 == EntId[3:0] ? dataArray_10_6_cachedata_MPORT_data : _GEN_1461; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1463 = _GEN_1872 & 4'h7 == EntId[3:0] ? dataArray_10_7_cachedata_MPORT_data : _GEN_1462; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1464 = _GEN_1872 & 4'h8 == EntId[3:0] ? dataArray_10_8_cachedata_MPORT_data : _GEN_1463; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1465 = _GEN_1872 & 4'h9 == EntId[3:0] ? dataArray_10_9_cachedata_MPORT_data : _GEN_1464; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1466 = _GEN_1872 & 4'ha == EntId[3:0] ? dataArray_10_10_cachedata_MPORT_data : _GEN_1465; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1467 = _GEN_1872 & 4'hb == EntId[3:0] ? dataArray_10_11_cachedata_MPORT_data : _GEN_1466; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1468 = _GEN_1872 & 4'hc == EntId[3:0] ? dataArray_10_12_cachedata_MPORT_data : _GEN_1467; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1469 = _GEN_1872 & 4'hd == EntId[3:0] ? dataArray_10_13_cachedata_MPORT_data : _GEN_1468; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1470 = _GEN_1872 & 4'he == EntId[3:0] ? dataArray_10_14_cachedata_MPORT_data : _GEN_1469; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1471 = _GEN_1872 & 4'hf == EntId[3:0] ? dataArray_10_15_cachedata_MPORT_data : _GEN_1470; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1472 = _GEN_1904 & 4'h0 == EntId[3:0] ? dataArray_11_0_cachedata_MPORT_data : _GEN_1471; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1473 = _GEN_1904 & 4'h1 == EntId[3:0] ? dataArray_11_1_cachedata_MPORT_data : _GEN_1472; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1474 = _GEN_1904 & 4'h2 == EntId[3:0] ? dataArray_11_2_cachedata_MPORT_data : _GEN_1473; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1475 = _GEN_1904 & 4'h3 == EntId[3:0] ? dataArray_11_3_cachedata_MPORT_data : _GEN_1474; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1476 = _GEN_1904 & 4'h4 == EntId[3:0] ? dataArray_11_4_cachedata_MPORT_data : _GEN_1475; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1477 = _GEN_1904 & 4'h5 == EntId[3:0] ? dataArray_11_5_cachedata_MPORT_data : _GEN_1476; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1478 = _GEN_1904 & 4'h6 == EntId[3:0] ? dataArray_11_6_cachedata_MPORT_data : _GEN_1477; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1479 = _GEN_1904 & 4'h7 == EntId[3:0] ? dataArray_11_7_cachedata_MPORT_data : _GEN_1478; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1480 = _GEN_1904 & 4'h8 == EntId[3:0] ? dataArray_11_8_cachedata_MPORT_data : _GEN_1479; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1481 = _GEN_1904 & 4'h9 == EntId[3:0] ? dataArray_11_9_cachedata_MPORT_data : _GEN_1480; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1482 = _GEN_1904 & 4'ha == EntId[3:0] ? dataArray_11_10_cachedata_MPORT_data : _GEN_1481; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1483 = _GEN_1904 & 4'hb == EntId[3:0] ? dataArray_11_11_cachedata_MPORT_data : _GEN_1482; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1484 = _GEN_1904 & 4'hc == EntId[3:0] ? dataArray_11_12_cachedata_MPORT_data : _GEN_1483; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1485 = _GEN_1904 & 4'hd == EntId[3:0] ? dataArray_11_13_cachedata_MPORT_data : _GEN_1484; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1486 = _GEN_1904 & 4'he == EntId[3:0] ? dataArray_11_14_cachedata_MPORT_data : _GEN_1485; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1487 = _GEN_1904 & 4'hf == EntId[3:0] ? dataArray_11_15_cachedata_MPORT_data : _GEN_1486; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1488 = _GEN_1936 & 4'h0 == EntId[3:0] ? dataArray_12_0_cachedata_MPORT_data : _GEN_1487; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1489 = _GEN_1936 & 4'h1 == EntId[3:0] ? dataArray_12_1_cachedata_MPORT_data : _GEN_1488; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1490 = _GEN_1936 & 4'h2 == EntId[3:0] ? dataArray_12_2_cachedata_MPORT_data : _GEN_1489; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1491 = _GEN_1936 & 4'h3 == EntId[3:0] ? dataArray_12_3_cachedata_MPORT_data : _GEN_1490; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1492 = _GEN_1936 & 4'h4 == EntId[3:0] ? dataArray_12_4_cachedata_MPORT_data : _GEN_1491; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1493 = _GEN_1936 & 4'h5 == EntId[3:0] ? dataArray_12_5_cachedata_MPORT_data : _GEN_1492; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1494 = _GEN_1936 & 4'h6 == EntId[3:0] ? dataArray_12_6_cachedata_MPORT_data : _GEN_1493; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1495 = _GEN_1936 & 4'h7 == EntId[3:0] ? dataArray_12_7_cachedata_MPORT_data : _GEN_1494; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1496 = _GEN_1936 & 4'h8 == EntId[3:0] ? dataArray_12_8_cachedata_MPORT_data : _GEN_1495; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1497 = _GEN_1936 & 4'h9 == EntId[3:0] ? dataArray_12_9_cachedata_MPORT_data : _GEN_1496; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1498 = _GEN_1936 & 4'ha == EntId[3:0] ? dataArray_12_10_cachedata_MPORT_data : _GEN_1497; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1499 = _GEN_1936 & 4'hb == EntId[3:0] ? dataArray_12_11_cachedata_MPORT_data : _GEN_1498; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1500 = _GEN_1936 & 4'hc == EntId[3:0] ? dataArray_12_12_cachedata_MPORT_data : _GEN_1499; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1501 = _GEN_1936 & 4'hd == EntId[3:0] ? dataArray_12_13_cachedata_MPORT_data : _GEN_1500; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1502 = _GEN_1936 & 4'he == EntId[3:0] ? dataArray_12_14_cachedata_MPORT_data : _GEN_1501; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1503 = _GEN_1936 & 4'hf == EntId[3:0] ? dataArray_12_15_cachedata_MPORT_data : _GEN_1502; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1504 = _GEN_1968 & 4'h0 == EntId[3:0] ? dataArray_13_0_cachedata_MPORT_data : _GEN_1503; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1505 = _GEN_1968 & 4'h1 == EntId[3:0] ? dataArray_13_1_cachedata_MPORT_data : _GEN_1504; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1506 = _GEN_1968 & 4'h2 == EntId[3:0] ? dataArray_13_2_cachedata_MPORT_data : _GEN_1505; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1507 = _GEN_1968 & 4'h3 == EntId[3:0] ? dataArray_13_3_cachedata_MPORT_data : _GEN_1506; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1508 = _GEN_1968 & 4'h4 == EntId[3:0] ? dataArray_13_4_cachedata_MPORT_data : _GEN_1507; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1509 = _GEN_1968 & 4'h5 == EntId[3:0] ? dataArray_13_5_cachedata_MPORT_data : _GEN_1508; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1510 = _GEN_1968 & 4'h6 == EntId[3:0] ? dataArray_13_6_cachedata_MPORT_data : _GEN_1509; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1511 = _GEN_1968 & 4'h7 == EntId[3:0] ? dataArray_13_7_cachedata_MPORT_data : _GEN_1510; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1512 = _GEN_1968 & 4'h8 == EntId[3:0] ? dataArray_13_8_cachedata_MPORT_data : _GEN_1511; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1513 = _GEN_1968 & 4'h9 == EntId[3:0] ? dataArray_13_9_cachedata_MPORT_data : _GEN_1512; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1514 = _GEN_1968 & 4'ha == EntId[3:0] ? dataArray_13_10_cachedata_MPORT_data : _GEN_1513; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1515 = _GEN_1968 & 4'hb == EntId[3:0] ? dataArray_13_11_cachedata_MPORT_data : _GEN_1514; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1516 = _GEN_1968 & 4'hc == EntId[3:0] ? dataArray_13_12_cachedata_MPORT_data : _GEN_1515; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1517 = _GEN_1968 & 4'hd == EntId[3:0] ? dataArray_13_13_cachedata_MPORT_data : _GEN_1516; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1518 = _GEN_1968 & 4'he == EntId[3:0] ? dataArray_13_14_cachedata_MPORT_data : _GEN_1517; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1519 = _GEN_1968 & 4'hf == EntId[3:0] ? dataArray_13_15_cachedata_MPORT_data : _GEN_1518; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1520 = _GEN_2000 & 4'h0 == EntId[3:0] ? dataArray_14_0_cachedata_MPORT_data : _GEN_1519; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1521 = _GEN_2000 & 4'h1 == EntId[3:0] ? dataArray_14_1_cachedata_MPORT_data : _GEN_1520; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1522 = _GEN_2000 & 4'h2 == EntId[3:0] ? dataArray_14_2_cachedata_MPORT_data : _GEN_1521; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1523 = _GEN_2000 & 4'h3 == EntId[3:0] ? dataArray_14_3_cachedata_MPORT_data : _GEN_1522; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1524 = _GEN_2000 & 4'h4 == EntId[3:0] ? dataArray_14_4_cachedata_MPORT_data : _GEN_1523; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1525 = _GEN_2000 & 4'h5 == EntId[3:0] ? dataArray_14_5_cachedata_MPORT_data : _GEN_1524; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1526 = _GEN_2000 & 4'h6 == EntId[3:0] ? dataArray_14_6_cachedata_MPORT_data : _GEN_1525; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1527 = _GEN_2000 & 4'h7 == EntId[3:0] ? dataArray_14_7_cachedata_MPORT_data : _GEN_1526; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1528 = _GEN_2000 & 4'h8 == EntId[3:0] ? dataArray_14_8_cachedata_MPORT_data : _GEN_1527; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1529 = _GEN_2000 & 4'h9 == EntId[3:0] ? dataArray_14_9_cachedata_MPORT_data : _GEN_1528; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1530 = _GEN_2000 & 4'ha == EntId[3:0] ? dataArray_14_10_cachedata_MPORT_data : _GEN_1529; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1531 = _GEN_2000 & 4'hb == EntId[3:0] ? dataArray_14_11_cachedata_MPORT_data : _GEN_1530; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1532 = _GEN_2000 & 4'hc == EntId[3:0] ? dataArray_14_12_cachedata_MPORT_data : _GEN_1531; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1533 = _GEN_2000 & 4'hd == EntId[3:0] ? dataArray_14_13_cachedata_MPORT_data : _GEN_1532; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1534 = _GEN_2000 & 4'he == EntId[3:0] ? dataArray_14_14_cachedata_MPORT_data : _GEN_1533; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1535 = _GEN_2000 & 4'hf == EntId[3:0] ? dataArray_14_15_cachedata_MPORT_data : _GEN_1534; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1536 = _GEN_2032 & 4'h0 == EntId[3:0] ? dataArray_15_0_cachedata_MPORT_data : _GEN_1535; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1537 = _GEN_2032 & 4'h1 == EntId[3:0] ? dataArray_15_1_cachedata_MPORT_data : _GEN_1536; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1538 = _GEN_2032 & 4'h2 == EntId[3:0] ? dataArray_15_2_cachedata_MPORT_data : _GEN_1537; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1539 = _GEN_2032 & 4'h3 == EntId[3:0] ? dataArray_15_3_cachedata_MPORT_data : _GEN_1538; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1540 = _GEN_2032 & 4'h4 == EntId[3:0] ? dataArray_15_4_cachedata_MPORT_data : _GEN_1539; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1541 = _GEN_2032 & 4'h5 == EntId[3:0] ? dataArray_15_5_cachedata_MPORT_data : _GEN_1540; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1542 = _GEN_2032 & 4'h6 == EntId[3:0] ? dataArray_15_6_cachedata_MPORT_data : _GEN_1541; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1543 = _GEN_2032 & 4'h7 == EntId[3:0] ? dataArray_15_7_cachedata_MPORT_data : _GEN_1542; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1544 = _GEN_2032 & 4'h8 == EntId[3:0] ? dataArray_15_8_cachedata_MPORT_data : _GEN_1543; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1545 = _GEN_2032 & 4'h9 == EntId[3:0] ? dataArray_15_9_cachedata_MPORT_data : _GEN_1544; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1546 = _GEN_2032 & 4'ha == EntId[3:0] ? dataArray_15_10_cachedata_MPORT_data : _GEN_1545; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1547 = _GEN_2032 & 4'hb == EntId[3:0] ? dataArray_15_11_cachedata_MPORT_data : _GEN_1546; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1548 = _GEN_2032 & 4'hc == EntId[3:0] ? dataArray_15_12_cachedata_MPORT_data : _GEN_1547; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1549 = _GEN_2032 & 4'hd == EntId[3:0] ? dataArray_15_13_cachedata_MPORT_data : _GEN_1548; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1550 = _GEN_2032 & 4'he == EntId[3:0] ? dataArray_15_14_cachedata_MPORT_data : _GEN_1549; // @[cache.scala 108:{28,28}]
  wire [31:0] _GEN_1551 = _GEN_2032 & 4'hf == EntId[3:0] ? dataArray_15_15_cachedata_MPORT_data : _GEN_1550; // @[cache.scala 108:{28,28}]
  assign dataArray_0_0_cachedata_MPORT_en = dataArray_0_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_0_cachedata_MPORT_addr = dataArray_0_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_0_cachedata_MPORT_data = dataArray_0_0[dataArray_0_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_0_MPORT_addr = replace_set;
  assign dataArray_0_0_MPORT_mask = _GEN_1552 & _GEN_1553;
  assign dataArray_0_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_1_cachedata_MPORT_en = dataArray_0_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_1_cachedata_MPORT_addr = dataArray_0_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_1_cachedata_MPORT_data = dataArray_0_1[dataArray_0_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_1_MPORT_addr = replace_set;
  assign dataArray_0_1_MPORT_mask = _GEN_1552 & _GEN_1555;
  assign dataArray_0_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_2_cachedata_MPORT_en = dataArray_0_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_2_cachedata_MPORT_addr = dataArray_0_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_2_cachedata_MPORT_data = dataArray_0_2[dataArray_0_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_2_MPORT_addr = replace_set;
  assign dataArray_0_2_MPORT_mask = _GEN_1552 & _GEN_1557;
  assign dataArray_0_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_3_cachedata_MPORT_en = dataArray_0_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_3_cachedata_MPORT_addr = dataArray_0_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_3_cachedata_MPORT_data = dataArray_0_3[dataArray_0_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_3_MPORT_addr = replace_set;
  assign dataArray_0_3_MPORT_mask = _GEN_1552 & _GEN_1559;
  assign dataArray_0_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_4_cachedata_MPORT_en = dataArray_0_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_4_cachedata_MPORT_addr = dataArray_0_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_4_cachedata_MPORT_data = dataArray_0_4[dataArray_0_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_4_MPORT_addr = replace_set;
  assign dataArray_0_4_MPORT_mask = _GEN_1552 & _GEN_1561;
  assign dataArray_0_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_5_cachedata_MPORT_en = dataArray_0_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_5_cachedata_MPORT_addr = dataArray_0_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_5_cachedata_MPORT_data = dataArray_0_5[dataArray_0_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_5_MPORT_addr = replace_set;
  assign dataArray_0_5_MPORT_mask = _GEN_1552 & _GEN_1563;
  assign dataArray_0_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_6_cachedata_MPORT_en = dataArray_0_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_6_cachedata_MPORT_addr = dataArray_0_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_6_cachedata_MPORT_data = dataArray_0_6[dataArray_0_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_6_MPORT_addr = replace_set;
  assign dataArray_0_6_MPORT_mask = _GEN_1552 & _GEN_1565;
  assign dataArray_0_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_7_cachedata_MPORT_en = dataArray_0_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_7_cachedata_MPORT_addr = dataArray_0_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_7_cachedata_MPORT_data = dataArray_0_7[dataArray_0_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_7_MPORT_addr = replace_set;
  assign dataArray_0_7_MPORT_mask = _GEN_1552 & _GEN_1567;
  assign dataArray_0_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_8_cachedata_MPORT_en = dataArray_0_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_8_cachedata_MPORT_addr = dataArray_0_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_8_cachedata_MPORT_data = dataArray_0_8[dataArray_0_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_8_MPORT_addr = replace_set;
  assign dataArray_0_8_MPORT_mask = _GEN_1552 & _GEN_1569;
  assign dataArray_0_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_9_cachedata_MPORT_en = dataArray_0_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_9_cachedata_MPORT_addr = dataArray_0_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_9_cachedata_MPORT_data = dataArray_0_9[dataArray_0_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_9_MPORT_addr = replace_set;
  assign dataArray_0_9_MPORT_mask = _GEN_1552 & _GEN_1571;
  assign dataArray_0_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_10_cachedata_MPORT_en = dataArray_0_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_10_cachedata_MPORT_addr = dataArray_0_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_10_cachedata_MPORT_data = dataArray_0_10[dataArray_0_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_10_MPORT_addr = replace_set;
  assign dataArray_0_10_MPORT_mask = _GEN_1552 & _GEN_1573;
  assign dataArray_0_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_11_cachedata_MPORT_en = dataArray_0_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_11_cachedata_MPORT_addr = dataArray_0_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_11_cachedata_MPORT_data = dataArray_0_11[dataArray_0_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_11_MPORT_addr = replace_set;
  assign dataArray_0_11_MPORT_mask = _GEN_1552 & _GEN_1575;
  assign dataArray_0_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_12_cachedata_MPORT_en = dataArray_0_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_12_cachedata_MPORT_addr = dataArray_0_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_12_cachedata_MPORT_data = dataArray_0_12[dataArray_0_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_12_MPORT_addr = replace_set;
  assign dataArray_0_12_MPORT_mask = _GEN_1552 & _GEN_1577;
  assign dataArray_0_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_13_cachedata_MPORT_en = dataArray_0_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_13_cachedata_MPORT_addr = dataArray_0_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_13_cachedata_MPORT_data = dataArray_0_13[dataArray_0_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_13_MPORT_addr = replace_set;
  assign dataArray_0_13_MPORT_mask = _GEN_1552 & _GEN_1579;
  assign dataArray_0_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_14_cachedata_MPORT_en = dataArray_0_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_14_cachedata_MPORT_addr = dataArray_0_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_14_cachedata_MPORT_data = dataArray_0_14[dataArray_0_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_14_MPORT_addr = replace_set;
  assign dataArray_0_14_MPORT_mask = _GEN_1552 & _GEN_1581;
  assign dataArray_0_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_0_15_cachedata_MPORT_en = dataArray_0_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_0_15_cachedata_MPORT_addr = dataArray_0_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_0_15_cachedata_MPORT_data = dataArray_0_15[dataArray_0_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_0_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_0_15_MPORT_addr = replace_set;
  assign dataArray_0_15_MPORT_mask = _GEN_1552 & _GEN_1583;
  assign dataArray_0_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_0_cachedata_MPORT_en = dataArray_1_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_0_cachedata_MPORT_addr = dataArray_1_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_0_cachedata_MPORT_data = dataArray_1_0[dataArray_1_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_0_MPORT_addr = replace_set;
  assign dataArray_1_0_MPORT_mask = _GEN_1584 & _GEN_1553;
  assign dataArray_1_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_1_cachedata_MPORT_en = dataArray_1_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_1_cachedata_MPORT_addr = dataArray_1_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_1_cachedata_MPORT_data = dataArray_1_1[dataArray_1_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_1_MPORT_addr = replace_set;
  assign dataArray_1_1_MPORT_mask = _GEN_1584 & _GEN_1555;
  assign dataArray_1_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_2_cachedata_MPORT_en = dataArray_1_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_2_cachedata_MPORT_addr = dataArray_1_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_2_cachedata_MPORT_data = dataArray_1_2[dataArray_1_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_2_MPORT_addr = replace_set;
  assign dataArray_1_2_MPORT_mask = _GEN_1584 & _GEN_1557;
  assign dataArray_1_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_3_cachedata_MPORT_en = dataArray_1_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_3_cachedata_MPORT_addr = dataArray_1_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_3_cachedata_MPORT_data = dataArray_1_3[dataArray_1_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_3_MPORT_addr = replace_set;
  assign dataArray_1_3_MPORT_mask = _GEN_1584 & _GEN_1559;
  assign dataArray_1_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_4_cachedata_MPORT_en = dataArray_1_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_4_cachedata_MPORT_addr = dataArray_1_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_4_cachedata_MPORT_data = dataArray_1_4[dataArray_1_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_4_MPORT_addr = replace_set;
  assign dataArray_1_4_MPORT_mask = _GEN_1584 & _GEN_1561;
  assign dataArray_1_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_5_cachedata_MPORT_en = dataArray_1_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_5_cachedata_MPORT_addr = dataArray_1_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_5_cachedata_MPORT_data = dataArray_1_5[dataArray_1_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_5_MPORT_addr = replace_set;
  assign dataArray_1_5_MPORT_mask = _GEN_1584 & _GEN_1563;
  assign dataArray_1_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_6_cachedata_MPORT_en = dataArray_1_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_6_cachedata_MPORT_addr = dataArray_1_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_6_cachedata_MPORT_data = dataArray_1_6[dataArray_1_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_6_MPORT_addr = replace_set;
  assign dataArray_1_6_MPORT_mask = _GEN_1584 & _GEN_1565;
  assign dataArray_1_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_7_cachedata_MPORT_en = dataArray_1_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_7_cachedata_MPORT_addr = dataArray_1_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_7_cachedata_MPORT_data = dataArray_1_7[dataArray_1_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_7_MPORT_addr = replace_set;
  assign dataArray_1_7_MPORT_mask = _GEN_1584 & _GEN_1567;
  assign dataArray_1_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_8_cachedata_MPORT_en = dataArray_1_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_8_cachedata_MPORT_addr = dataArray_1_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_8_cachedata_MPORT_data = dataArray_1_8[dataArray_1_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_8_MPORT_addr = replace_set;
  assign dataArray_1_8_MPORT_mask = _GEN_1584 & _GEN_1569;
  assign dataArray_1_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_9_cachedata_MPORT_en = dataArray_1_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_9_cachedata_MPORT_addr = dataArray_1_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_9_cachedata_MPORT_data = dataArray_1_9[dataArray_1_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_9_MPORT_addr = replace_set;
  assign dataArray_1_9_MPORT_mask = _GEN_1584 & _GEN_1571;
  assign dataArray_1_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_10_cachedata_MPORT_en = dataArray_1_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_10_cachedata_MPORT_addr = dataArray_1_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_10_cachedata_MPORT_data = dataArray_1_10[dataArray_1_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_10_MPORT_addr = replace_set;
  assign dataArray_1_10_MPORT_mask = _GEN_1584 & _GEN_1573;
  assign dataArray_1_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_11_cachedata_MPORT_en = dataArray_1_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_11_cachedata_MPORT_addr = dataArray_1_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_11_cachedata_MPORT_data = dataArray_1_11[dataArray_1_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_11_MPORT_addr = replace_set;
  assign dataArray_1_11_MPORT_mask = _GEN_1584 & _GEN_1575;
  assign dataArray_1_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_12_cachedata_MPORT_en = dataArray_1_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_12_cachedata_MPORT_addr = dataArray_1_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_12_cachedata_MPORT_data = dataArray_1_12[dataArray_1_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_12_MPORT_addr = replace_set;
  assign dataArray_1_12_MPORT_mask = _GEN_1584 & _GEN_1577;
  assign dataArray_1_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_13_cachedata_MPORT_en = dataArray_1_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_13_cachedata_MPORT_addr = dataArray_1_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_13_cachedata_MPORT_data = dataArray_1_13[dataArray_1_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_13_MPORT_addr = replace_set;
  assign dataArray_1_13_MPORT_mask = _GEN_1584 & _GEN_1579;
  assign dataArray_1_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_14_cachedata_MPORT_en = dataArray_1_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_14_cachedata_MPORT_addr = dataArray_1_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_14_cachedata_MPORT_data = dataArray_1_14[dataArray_1_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_14_MPORT_addr = replace_set;
  assign dataArray_1_14_MPORT_mask = _GEN_1584 & _GEN_1581;
  assign dataArray_1_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_1_15_cachedata_MPORT_en = dataArray_1_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_1_15_cachedata_MPORT_addr = dataArray_1_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_1_15_cachedata_MPORT_data = dataArray_1_15[dataArray_1_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_1_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_1_15_MPORT_addr = replace_set;
  assign dataArray_1_15_MPORT_mask = _GEN_1584 & _GEN_1583;
  assign dataArray_1_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_0_cachedata_MPORT_en = dataArray_2_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_0_cachedata_MPORT_addr = dataArray_2_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_0_cachedata_MPORT_data = dataArray_2_0[dataArray_2_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_0_MPORT_addr = replace_set;
  assign dataArray_2_0_MPORT_mask = _GEN_1616 & _GEN_1553;
  assign dataArray_2_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_1_cachedata_MPORT_en = dataArray_2_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_1_cachedata_MPORT_addr = dataArray_2_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_1_cachedata_MPORT_data = dataArray_2_1[dataArray_2_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_1_MPORT_addr = replace_set;
  assign dataArray_2_1_MPORT_mask = _GEN_1616 & _GEN_1555;
  assign dataArray_2_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_2_cachedata_MPORT_en = dataArray_2_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_2_cachedata_MPORT_addr = dataArray_2_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_2_cachedata_MPORT_data = dataArray_2_2[dataArray_2_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_2_MPORT_addr = replace_set;
  assign dataArray_2_2_MPORT_mask = _GEN_1616 & _GEN_1557;
  assign dataArray_2_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_3_cachedata_MPORT_en = dataArray_2_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_3_cachedata_MPORT_addr = dataArray_2_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_3_cachedata_MPORT_data = dataArray_2_3[dataArray_2_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_3_MPORT_addr = replace_set;
  assign dataArray_2_3_MPORT_mask = _GEN_1616 & _GEN_1559;
  assign dataArray_2_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_4_cachedata_MPORT_en = dataArray_2_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_4_cachedata_MPORT_addr = dataArray_2_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_4_cachedata_MPORT_data = dataArray_2_4[dataArray_2_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_4_MPORT_addr = replace_set;
  assign dataArray_2_4_MPORT_mask = _GEN_1616 & _GEN_1561;
  assign dataArray_2_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_5_cachedata_MPORT_en = dataArray_2_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_5_cachedata_MPORT_addr = dataArray_2_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_5_cachedata_MPORT_data = dataArray_2_5[dataArray_2_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_5_MPORT_addr = replace_set;
  assign dataArray_2_5_MPORT_mask = _GEN_1616 & _GEN_1563;
  assign dataArray_2_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_6_cachedata_MPORT_en = dataArray_2_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_6_cachedata_MPORT_addr = dataArray_2_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_6_cachedata_MPORT_data = dataArray_2_6[dataArray_2_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_6_MPORT_addr = replace_set;
  assign dataArray_2_6_MPORT_mask = _GEN_1616 & _GEN_1565;
  assign dataArray_2_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_7_cachedata_MPORT_en = dataArray_2_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_7_cachedata_MPORT_addr = dataArray_2_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_7_cachedata_MPORT_data = dataArray_2_7[dataArray_2_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_7_MPORT_addr = replace_set;
  assign dataArray_2_7_MPORT_mask = _GEN_1616 & _GEN_1567;
  assign dataArray_2_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_8_cachedata_MPORT_en = dataArray_2_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_8_cachedata_MPORT_addr = dataArray_2_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_8_cachedata_MPORT_data = dataArray_2_8[dataArray_2_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_8_MPORT_addr = replace_set;
  assign dataArray_2_8_MPORT_mask = _GEN_1616 & _GEN_1569;
  assign dataArray_2_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_9_cachedata_MPORT_en = dataArray_2_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_9_cachedata_MPORT_addr = dataArray_2_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_9_cachedata_MPORT_data = dataArray_2_9[dataArray_2_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_9_MPORT_addr = replace_set;
  assign dataArray_2_9_MPORT_mask = _GEN_1616 & _GEN_1571;
  assign dataArray_2_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_10_cachedata_MPORT_en = dataArray_2_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_10_cachedata_MPORT_addr = dataArray_2_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_10_cachedata_MPORT_data = dataArray_2_10[dataArray_2_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_10_MPORT_addr = replace_set;
  assign dataArray_2_10_MPORT_mask = _GEN_1616 & _GEN_1573;
  assign dataArray_2_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_11_cachedata_MPORT_en = dataArray_2_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_11_cachedata_MPORT_addr = dataArray_2_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_11_cachedata_MPORT_data = dataArray_2_11[dataArray_2_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_11_MPORT_addr = replace_set;
  assign dataArray_2_11_MPORT_mask = _GEN_1616 & _GEN_1575;
  assign dataArray_2_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_12_cachedata_MPORT_en = dataArray_2_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_12_cachedata_MPORT_addr = dataArray_2_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_12_cachedata_MPORT_data = dataArray_2_12[dataArray_2_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_12_MPORT_addr = replace_set;
  assign dataArray_2_12_MPORT_mask = _GEN_1616 & _GEN_1577;
  assign dataArray_2_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_13_cachedata_MPORT_en = dataArray_2_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_13_cachedata_MPORT_addr = dataArray_2_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_13_cachedata_MPORT_data = dataArray_2_13[dataArray_2_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_13_MPORT_addr = replace_set;
  assign dataArray_2_13_MPORT_mask = _GEN_1616 & _GEN_1579;
  assign dataArray_2_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_14_cachedata_MPORT_en = dataArray_2_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_14_cachedata_MPORT_addr = dataArray_2_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_14_cachedata_MPORT_data = dataArray_2_14[dataArray_2_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_14_MPORT_addr = replace_set;
  assign dataArray_2_14_MPORT_mask = _GEN_1616 & _GEN_1581;
  assign dataArray_2_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_2_15_cachedata_MPORT_en = dataArray_2_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_2_15_cachedata_MPORT_addr = dataArray_2_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_2_15_cachedata_MPORT_data = dataArray_2_15[dataArray_2_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_2_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_2_15_MPORT_addr = replace_set;
  assign dataArray_2_15_MPORT_mask = _GEN_1616 & _GEN_1583;
  assign dataArray_2_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_0_cachedata_MPORT_en = dataArray_3_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_0_cachedata_MPORT_addr = dataArray_3_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_0_cachedata_MPORT_data = dataArray_3_0[dataArray_3_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_0_MPORT_addr = replace_set;
  assign dataArray_3_0_MPORT_mask = _GEN_1648 & _GEN_1553;
  assign dataArray_3_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_1_cachedata_MPORT_en = dataArray_3_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_1_cachedata_MPORT_addr = dataArray_3_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_1_cachedata_MPORT_data = dataArray_3_1[dataArray_3_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_1_MPORT_addr = replace_set;
  assign dataArray_3_1_MPORT_mask = _GEN_1648 & _GEN_1555;
  assign dataArray_3_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_2_cachedata_MPORT_en = dataArray_3_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_2_cachedata_MPORT_addr = dataArray_3_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_2_cachedata_MPORT_data = dataArray_3_2[dataArray_3_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_2_MPORT_addr = replace_set;
  assign dataArray_3_2_MPORT_mask = _GEN_1648 & _GEN_1557;
  assign dataArray_3_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_3_cachedata_MPORT_en = dataArray_3_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_3_cachedata_MPORT_addr = dataArray_3_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_3_cachedata_MPORT_data = dataArray_3_3[dataArray_3_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_3_MPORT_addr = replace_set;
  assign dataArray_3_3_MPORT_mask = _GEN_1648 & _GEN_1559;
  assign dataArray_3_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_4_cachedata_MPORT_en = dataArray_3_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_4_cachedata_MPORT_addr = dataArray_3_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_4_cachedata_MPORT_data = dataArray_3_4[dataArray_3_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_4_MPORT_addr = replace_set;
  assign dataArray_3_4_MPORT_mask = _GEN_1648 & _GEN_1561;
  assign dataArray_3_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_5_cachedata_MPORT_en = dataArray_3_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_5_cachedata_MPORT_addr = dataArray_3_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_5_cachedata_MPORT_data = dataArray_3_5[dataArray_3_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_5_MPORT_addr = replace_set;
  assign dataArray_3_5_MPORT_mask = _GEN_1648 & _GEN_1563;
  assign dataArray_3_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_6_cachedata_MPORT_en = dataArray_3_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_6_cachedata_MPORT_addr = dataArray_3_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_6_cachedata_MPORT_data = dataArray_3_6[dataArray_3_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_6_MPORT_addr = replace_set;
  assign dataArray_3_6_MPORT_mask = _GEN_1648 & _GEN_1565;
  assign dataArray_3_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_7_cachedata_MPORT_en = dataArray_3_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_7_cachedata_MPORT_addr = dataArray_3_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_7_cachedata_MPORT_data = dataArray_3_7[dataArray_3_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_7_MPORT_addr = replace_set;
  assign dataArray_3_7_MPORT_mask = _GEN_1648 & _GEN_1567;
  assign dataArray_3_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_8_cachedata_MPORT_en = dataArray_3_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_8_cachedata_MPORT_addr = dataArray_3_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_8_cachedata_MPORT_data = dataArray_3_8[dataArray_3_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_8_MPORT_addr = replace_set;
  assign dataArray_3_8_MPORT_mask = _GEN_1648 & _GEN_1569;
  assign dataArray_3_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_9_cachedata_MPORT_en = dataArray_3_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_9_cachedata_MPORT_addr = dataArray_3_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_9_cachedata_MPORT_data = dataArray_3_9[dataArray_3_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_9_MPORT_addr = replace_set;
  assign dataArray_3_9_MPORT_mask = _GEN_1648 & _GEN_1571;
  assign dataArray_3_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_10_cachedata_MPORT_en = dataArray_3_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_10_cachedata_MPORT_addr = dataArray_3_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_10_cachedata_MPORT_data = dataArray_3_10[dataArray_3_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_10_MPORT_addr = replace_set;
  assign dataArray_3_10_MPORT_mask = _GEN_1648 & _GEN_1573;
  assign dataArray_3_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_11_cachedata_MPORT_en = dataArray_3_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_11_cachedata_MPORT_addr = dataArray_3_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_11_cachedata_MPORT_data = dataArray_3_11[dataArray_3_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_11_MPORT_addr = replace_set;
  assign dataArray_3_11_MPORT_mask = _GEN_1648 & _GEN_1575;
  assign dataArray_3_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_12_cachedata_MPORT_en = dataArray_3_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_12_cachedata_MPORT_addr = dataArray_3_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_12_cachedata_MPORT_data = dataArray_3_12[dataArray_3_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_12_MPORT_addr = replace_set;
  assign dataArray_3_12_MPORT_mask = _GEN_1648 & _GEN_1577;
  assign dataArray_3_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_13_cachedata_MPORT_en = dataArray_3_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_13_cachedata_MPORT_addr = dataArray_3_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_13_cachedata_MPORT_data = dataArray_3_13[dataArray_3_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_13_MPORT_addr = replace_set;
  assign dataArray_3_13_MPORT_mask = _GEN_1648 & _GEN_1579;
  assign dataArray_3_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_14_cachedata_MPORT_en = dataArray_3_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_14_cachedata_MPORT_addr = dataArray_3_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_14_cachedata_MPORT_data = dataArray_3_14[dataArray_3_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_14_MPORT_addr = replace_set;
  assign dataArray_3_14_MPORT_mask = _GEN_1648 & _GEN_1581;
  assign dataArray_3_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_3_15_cachedata_MPORT_en = dataArray_3_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_3_15_cachedata_MPORT_addr = dataArray_3_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_3_15_cachedata_MPORT_data = dataArray_3_15[dataArray_3_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_3_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_3_15_MPORT_addr = replace_set;
  assign dataArray_3_15_MPORT_mask = _GEN_1648 & _GEN_1583;
  assign dataArray_3_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_0_cachedata_MPORT_en = dataArray_4_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_0_cachedata_MPORT_addr = dataArray_4_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_0_cachedata_MPORT_data = dataArray_4_0[dataArray_4_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_0_MPORT_addr = replace_set;
  assign dataArray_4_0_MPORT_mask = _GEN_1680 & _GEN_1553;
  assign dataArray_4_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_1_cachedata_MPORT_en = dataArray_4_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_1_cachedata_MPORT_addr = dataArray_4_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_1_cachedata_MPORT_data = dataArray_4_1[dataArray_4_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_1_MPORT_addr = replace_set;
  assign dataArray_4_1_MPORT_mask = _GEN_1680 & _GEN_1555;
  assign dataArray_4_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_2_cachedata_MPORT_en = dataArray_4_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_2_cachedata_MPORT_addr = dataArray_4_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_2_cachedata_MPORT_data = dataArray_4_2[dataArray_4_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_2_MPORT_addr = replace_set;
  assign dataArray_4_2_MPORT_mask = _GEN_1680 & _GEN_1557;
  assign dataArray_4_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_3_cachedata_MPORT_en = dataArray_4_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_3_cachedata_MPORT_addr = dataArray_4_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_3_cachedata_MPORT_data = dataArray_4_3[dataArray_4_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_3_MPORT_addr = replace_set;
  assign dataArray_4_3_MPORT_mask = _GEN_1680 & _GEN_1559;
  assign dataArray_4_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_4_cachedata_MPORT_en = dataArray_4_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_4_cachedata_MPORT_addr = dataArray_4_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_4_cachedata_MPORT_data = dataArray_4_4[dataArray_4_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_4_MPORT_addr = replace_set;
  assign dataArray_4_4_MPORT_mask = _GEN_1680 & _GEN_1561;
  assign dataArray_4_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_5_cachedata_MPORT_en = dataArray_4_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_5_cachedata_MPORT_addr = dataArray_4_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_5_cachedata_MPORT_data = dataArray_4_5[dataArray_4_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_5_MPORT_addr = replace_set;
  assign dataArray_4_5_MPORT_mask = _GEN_1680 & _GEN_1563;
  assign dataArray_4_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_6_cachedata_MPORT_en = dataArray_4_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_6_cachedata_MPORT_addr = dataArray_4_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_6_cachedata_MPORT_data = dataArray_4_6[dataArray_4_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_6_MPORT_addr = replace_set;
  assign dataArray_4_6_MPORT_mask = _GEN_1680 & _GEN_1565;
  assign dataArray_4_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_7_cachedata_MPORT_en = dataArray_4_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_7_cachedata_MPORT_addr = dataArray_4_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_7_cachedata_MPORT_data = dataArray_4_7[dataArray_4_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_7_MPORT_addr = replace_set;
  assign dataArray_4_7_MPORT_mask = _GEN_1680 & _GEN_1567;
  assign dataArray_4_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_8_cachedata_MPORT_en = dataArray_4_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_8_cachedata_MPORT_addr = dataArray_4_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_8_cachedata_MPORT_data = dataArray_4_8[dataArray_4_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_8_MPORT_addr = replace_set;
  assign dataArray_4_8_MPORT_mask = _GEN_1680 & _GEN_1569;
  assign dataArray_4_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_9_cachedata_MPORT_en = dataArray_4_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_9_cachedata_MPORT_addr = dataArray_4_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_9_cachedata_MPORT_data = dataArray_4_9[dataArray_4_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_9_MPORT_addr = replace_set;
  assign dataArray_4_9_MPORT_mask = _GEN_1680 & _GEN_1571;
  assign dataArray_4_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_10_cachedata_MPORT_en = dataArray_4_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_10_cachedata_MPORT_addr = dataArray_4_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_10_cachedata_MPORT_data = dataArray_4_10[dataArray_4_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_10_MPORT_addr = replace_set;
  assign dataArray_4_10_MPORT_mask = _GEN_1680 & _GEN_1573;
  assign dataArray_4_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_11_cachedata_MPORT_en = dataArray_4_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_11_cachedata_MPORT_addr = dataArray_4_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_11_cachedata_MPORT_data = dataArray_4_11[dataArray_4_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_11_MPORT_addr = replace_set;
  assign dataArray_4_11_MPORT_mask = _GEN_1680 & _GEN_1575;
  assign dataArray_4_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_12_cachedata_MPORT_en = dataArray_4_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_12_cachedata_MPORT_addr = dataArray_4_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_12_cachedata_MPORT_data = dataArray_4_12[dataArray_4_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_12_MPORT_addr = replace_set;
  assign dataArray_4_12_MPORT_mask = _GEN_1680 & _GEN_1577;
  assign dataArray_4_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_13_cachedata_MPORT_en = dataArray_4_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_13_cachedata_MPORT_addr = dataArray_4_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_13_cachedata_MPORT_data = dataArray_4_13[dataArray_4_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_13_MPORT_addr = replace_set;
  assign dataArray_4_13_MPORT_mask = _GEN_1680 & _GEN_1579;
  assign dataArray_4_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_14_cachedata_MPORT_en = dataArray_4_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_14_cachedata_MPORT_addr = dataArray_4_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_14_cachedata_MPORT_data = dataArray_4_14[dataArray_4_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_14_MPORT_addr = replace_set;
  assign dataArray_4_14_MPORT_mask = _GEN_1680 & _GEN_1581;
  assign dataArray_4_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_4_15_cachedata_MPORT_en = dataArray_4_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_4_15_cachedata_MPORT_addr = dataArray_4_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_4_15_cachedata_MPORT_data = dataArray_4_15[dataArray_4_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_4_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_4_15_MPORT_addr = replace_set;
  assign dataArray_4_15_MPORT_mask = _GEN_1680 & _GEN_1583;
  assign dataArray_4_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_0_cachedata_MPORT_en = dataArray_5_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_0_cachedata_MPORT_addr = dataArray_5_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_0_cachedata_MPORT_data = dataArray_5_0[dataArray_5_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_0_MPORT_addr = replace_set;
  assign dataArray_5_0_MPORT_mask = _GEN_1712 & _GEN_1553;
  assign dataArray_5_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_1_cachedata_MPORT_en = dataArray_5_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_1_cachedata_MPORT_addr = dataArray_5_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_1_cachedata_MPORT_data = dataArray_5_1[dataArray_5_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_1_MPORT_addr = replace_set;
  assign dataArray_5_1_MPORT_mask = _GEN_1712 & _GEN_1555;
  assign dataArray_5_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_2_cachedata_MPORT_en = dataArray_5_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_2_cachedata_MPORT_addr = dataArray_5_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_2_cachedata_MPORT_data = dataArray_5_2[dataArray_5_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_2_MPORT_addr = replace_set;
  assign dataArray_5_2_MPORT_mask = _GEN_1712 & _GEN_1557;
  assign dataArray_5_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_3_cachedata_MPORT_en = dataArray_5_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_3_cachedata_MPORT_addr = dataArray_5_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_3_cachedata_MPORT_data = dataArray_5_3[dataArray_5_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_3_MPORT_addr = replace_set;
  assign dataArray_5_3_MPORT_mask = _GEN_1712 & _GEN_1559;
  assign dataArray_5_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_4_cachedata_MPORT_en = dataArray_5_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_4_cachedata_MPORT_addr = dataArray_5_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_4_cachedata_MPORT_data = dataArray_5_4[dataArray_5_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_4_MPORT_addr = replace_set;
  assign dataArray_5_4_MPORT_mask = _GEN_1712 & _GEN_1561;
  assign dataArray_5_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_5_cachedata_MPORT_en = dataArray_5_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_5_cachedata_MPORT_addr = dataArray_5_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_5_cachedata_MPORT_data = dataArray_5_5[dataArray_5_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_5_MPORT_addr = replace_set;
  assign dataArray_5_5_MPORT_mask = _GEN_1712 & _GEN_1563;
  assign dataArray_5_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_6_cachedata_MPORT_en = dataArray_5_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_6_cachedata_MPORT_addr = dataArray_5_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_6_cachedata_MPORT_data = dataArray_5_6[dataArray_5_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_6_MPORT_addr = replace_set;
  assign dataArray_5_6_MPORT_mask = _GEN_1712 & _GEN_1565;
  assign dataArray_5_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_7_cachedata_MPORT_en = dataArray_5_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_7_cachedata_MPORT_addr = dataArray_5_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_7_cachedata_MPORT_data = dataArray_5_7[dataArray_5_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_7_MPORT_addr = replace_set;
  assign dataArray_5_7_MPORT_mask = _GEN_1712 & _GEN_1567;
  assign dataArray_5_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_8_cachedata_MPORT_en = dataArray_5_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_8_cachedata_MPORT_addr = dataArray_5_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_8_cachedata_MPORT_data = dataArray_5_8[dataArray_5_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_8_MPORT_addr = replace_set;
  assign dataArray_5_8_MPORT_mask = _GEN_1712 & _GEN_1569;
  assign dataArray_5_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_9_cachedata_MPORT_en = dataArray_5_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_9_cachedata_MPORT_addr = dataArray_5_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_9_cachedata_MPORT_data = dataArray_5_9[dataArray_5_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_9_MPORT_addr = replace_set;
  assign dataArray_5_9_MPORT_mask = _GEN_1712 & _GEN_1571;
  assign dataArray_5_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_10_cachedata_MPORT_en = dataArray_5_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_10_cachedata_MPORT_addr = dataArray_5_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_10_cachedata_MPORT_data = dataArray_5_10[dataArray_5_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_10_MPORT_addr = replace_set;
  assign dataArray_5_10_MPORT_mask = _GEN_1712 & _GEN_1573;
  assign dataArray_5_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_11_cachedata_MPORT_en = dataArray_5_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_11_cachedata_MPORT_addr = dataArray_5_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_11_cachedata_MPORT_data = dataArray_5_11[dataArray_5_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_11_MPORT_addr = replace_set;
  assign dataArray_5_11_MPORT_mask = _GEN_1712 & _GEN_1575;
  assign dataArray_5_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_12_cachedata_MPORT_en = dataArray_5_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_12_cachedata_MPORT_addr = dataArray_5_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_12_cachedata_MPORT_data = dataArray_5_12[dataArray_5_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_12_MPORT_addr = replace_set;
  assign dataArray_5_12_MPORT_mask = _GEN_1712 & _GEN_1577;
  assign dataArray_5_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_13_cachedata_MPORT_en = dataArray_5_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_13_cachedata_MPORT_addr = dataArray_5_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_13_cachedata_MPORT_data = dataArray_5_13[dataArray_5_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_13_MPORT_addr = replace_set;
  assign dataArray_5_13_MPORT_mask = _GEN_1712 & _GEN_1579;
  assign dataArray_5_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_14_cachedata_MPORT_en = dataArray_5_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_14_cachedata_MPORT_addr = dataArray_5_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_14_cachedata_MPORT_data = dataArray_5_14[dataArray_5_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_14_MPORT_addr = replace_set;
  assign dataArray_5_14_MPORT_mask = _GEN_1712 & _GEN_1581;
  assign dataArray_5_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_5_15_cachedata_MPORT_en = dataArray_5_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_5_15_cachedata_MPORT_addr = dataArray_5_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_5_15_cachedata_MPORT_data = dataArray_5_15[dataArray_5_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_5_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_5_15_MPORT_addr = replace_set;
  assign dataArray_5_15_MPORT_mask = _GEN_1712 & _GEN_1583;
  assign dataArray_5_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_0_cachedata_MPORT_en = dataArray_6_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_0_cachedata_MPORT_addr = dataArray_6_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_0_cachedata_MPORT_data = dataArray_6_0[dataArray_6_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_0_MPORT_addr = replace_set;
  assign dataArray_6_0_MPORT_mask = _GEN_1744 & _GEN_1553;
  assign dataArray_6_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_1_cachedata_MPORT_en = dataArray_6_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_1_cachedata_MPORT_addr = dataArray_6_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_1_cachedata_MPORT_data = dataArray_6_1[dataArray_6_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_1_MPORT_addr = replace_set;
  assign dataArray_6_1_MPORT_mask = _GEN_1744 & _GEN_1555;
  assign dataArray_6_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_2_cachedata_MPORT_en = dataArray_6_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_2_cachedata_MPORT_addr = dataArray_6_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_2_cachedata_MPORT_data = dataArray_6_2[dataArray_6_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_2_MPORT_addr = replace_set;
  assign dataArray_6_2_MPORT_mask = _GEN_1744 & _GEN_1557;
  assign dataArray_6_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_3_cachedata_MPORT_en = dataArray_6_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_3_cachedata_MPORT_addr = dataArray_6_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_3_cachedata_MPORT_data = dataArray_6_3[dataArray_6_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_3_MPORT_addr = replace_set;
  assign dataArray_6_3_MPORT_mask = _GEN_1744 & _GEN_1559;
  assign dataArray_6_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_4_cachedata_MPORT_en = dataArray_6_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_4_cachedata_MPORT_addr = dataArray_6_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_4_cachedata_MPORT_data = dataArray_6_4[dataArray_6_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_4_MPORT_addr = replace_set;
  assign dataArray_6_4_MPORT_mask = _GEN_1744 & _GEN_1561;
  assign dataArray_6_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_5_cachedata_MPORT_en = dataArray_6_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_5_cachedata_MPORT_addr = dataArray_6_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_5_cachedata_MPORT_data = dataArray_6_5[dataArray_6_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_5_MPORT_addr = replace_set;
  assign dataArray_6_5_MPORT_mask = _GEN_1744 & _GEN_1563;
  assign dataArray_6_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_6_cachedata_MPORT_en = dataArray_6_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_6_cachedata_MPORT_addr = dataArray_6_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_6_cachedata_MPORT_data = dataArray_6_6[dataArray_6_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_6_MPORT_addr = replace_set;
  assign dataArray_6_6_MPORT_mask = _GEN_1744 & _GEN_1565;
  assign dataArray_6_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_7_cachedata_MPORT_en = dataArray_6_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_7_cachedata_MPORT_addr = dataArray_6_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_7_cachedata_MPORT_data = dataArray_6_7[dataArray_6_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_7_MPORT_addr = replace_set;
  assign dataArray_6_7_MPORT_mask = _GEN_1744 & _GEN_1567;
  assign dataArray_6_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_8_cachedata_MPORT_en = dataArray_6_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_8_cachedata_MPORT_addr = dataArray_6_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_8_cachedata_MPORT_data = dataArray_6_8[dataArray_6_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_8_MPORT_addr = replace_set;
  assign dataArray_6_8_MPORT_mask = _GEN_1744 & _GEN_1569;
  assign dataArray_6_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_9_cachedata_MPORT_en = dataArray_6_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_9_cachedata_MPORT_addr = dataArray_6_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_9_cachedata_MPORT_data = dataArray_6_9[dataArray_6_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_9_MPORT_addr = replace_set;
  assign dataArray_6_9_MPORT_mask = _GEN_1744 & _GEN_1571;
  assign dataArray_6_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_10_cachedata_MPORT_en = dataArray_6_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_10_cachedata_MPORT_addr = dataArray_6_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_10_cachedata_MPORT_data = dataArray_6_10[dataArray_6_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_10_MPORT_addr = replace_set;
  assign dataArray_6_10_MPORT_mask = _GEN_1744 & _GEN_1573;
  assign dataArray_6_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_11_cachedata_MPORT_en = dataArray_6_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_11_cachedata_MPORT_addr = dataArray_6_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_11_cachedata_MPORT_data = dataArray_6_11[dataArray_6_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_11_MPORT_addr = replace_set;
  assign dataArray_6_11_MPORT_mask = _GEN_1744 & _GEN_1575;
  assign dataArray_6_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_12_cachedata_MPORT_en = dataArray_6_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_12_cachedata_MPORT_addr = dataArray_6_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_12_cachedata_MPORT_data = dataArray_6_12[dataArray_6_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_12_MPORT_addr = replace_set;
  assign dataArray_6_12_MPORT_mask = _GEN_1744 & _GEN_1577;
  assign dataArray_6_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_13_cachedata_MPORT_en = dataArray_6_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_13_cachedata_MPORT_addr = dataArray_6_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_13_cachedata_MPORT_data = dataArray_6_13[dataArray_6_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_13_MPORT_addr = replace_set;
  assign dataArray_6_13_MPORT_mask = _GEN_1744 & _GEN_1579;
  assign dataArray_6_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_14_cachedata_MPORT_en = dataArray_6_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_14_cachedata_MPORT_addr = dataArray_6_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_14_cachedata_MPORT_data = dataArray_6_14[dataArray_6_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_14_MPORT_addr = replace_set;
  assign dataArray_6_14_MPORT_mask = _GEN_1744 & _GEN_1581;
  assign dataArray_6_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_6_15_cachedata_MPORT_en = dataArray_6_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_6_15_cachedata_MPORT_addr = dataArray_6_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_6_15_cachedata_MPORT_data = dataArray_6_15[dataArray_6_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_6_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_6_15_MPORT_addr = replace_set;
  assign dataArray_6_15_MPORT_mask = _GEN_1744 & _GEN_1583;
  assign dataArray_6_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_0_cachedata_MPORT_en = dataArray_7_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_0_cachedata_MPORT_addr = dataArray_7_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_0_cachedata_MPORT_data = dataArray_7_0[dataArray_7_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_0_MPORT_addr = replace_set;
  assign dataArray_7_0_MPORT_mask = _GEN_1776 & _GEN_1553;
  assign dataArray_7_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_1_cachedata_MPORT_en = dataArray_7_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_1_cachedata_MPORT_addr = dataArray_7_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_1_cachedata_MPORT_data = dataArray_7_1[dataArray_7_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_1_MPORT_addr = replace_set;
  assign dataArray_7_1_MPORT_mask = _GEN_1776 & _GEN_1555;
  assign dataArray_7_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_2_cachedata_MPORT_en = dataArray_7_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_2_cachedata_MPORT_addr = dataArray_7_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_2_cachedata_MPORT_data = dataArray_7_2[dataArray_7_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_2_MPORT_addr = replace_set;
  assign dataArray_7_2_MPORT_mask = _GEN_1776 & _GEN_1557;
  assign dataArray_7_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_3_cachedata_MPORT_en = dataArray_7_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_3_cachedata_MPORT_addr = dataArray_7_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_3_cachedata_MPORT_data = dataArray_7_3[dataArray_7_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_3_MPORT_addr = replace_set;
  assign dataArray_7_3_MPORT_mask = _GEN_1776 & _GEN_1559;
  assign dataArray_7_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_4_cachedata_MPORT_en = dataArray_7_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_4_cachedata_MPORT_addr = dataArray_7_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_4_cachedata_MPORT_data = dataArray_7_4[dataArray_7_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_4_MPORT_addr = replace_set;
  assign dataArray_7_4_MPORT_mask = _GEN_1776 & _GEN_1561;
  assign dataArray_7_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_5_cachedata_MPORT_en = dataArray_7_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_5_cachedata_MPORT_addr = dataArray_7_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_5_cachedata_MPORT_data = dataArray_7_5[dataArray_7_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_5_MPORT_addr = replace_set;
  assign dataArray_7_5_MPORT_mask = _GEN_1776 & _GEN_1563;
  assign dataArray_7_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_6_cachedata_MPORT_en = dataArray_7_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_6_cachedata_MPORT_addr = dataArray_7_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_6_cachedata_MPORT_data = dataArray_7_6[dataArray_7_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_6_MPORT_addr = replace_set;
  assign dataArray_7_6_MPORT_mask = _GEN_1776 & _GEN_1565;
  assign dataArray_7_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_7_cachedata_MPORT_en = dataArray_7_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_7_cachedata_MPORT_addr = dataArray_7_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_7_cachedata_MPORT_data = dataArray_7_7[dataArray_7_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_7_MPORT_addr = replace_set;
  assign dataArray_7_7_MPORT_mask = _GEN_1776 & _GEN_1567;
  assign dataArray_7_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_8_cachedata_MPORT_en = dataArray_7_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_8_cachedata_MPORT_addr = dataArray_7_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_8_cachedata_MPORT_data = dataArray_7_8[dataArray_7_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_8_MPORT_addr = replace_set;
  assign dataArray_7_8_MPORT_mask = _GEN_1776 & _GEN_1569;
  assign dataArray_7_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_9_cachedata_MPORT_en = dataArray_7_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_9_cachedata_MPORT_addr = dataArray_7_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_9_cachedata_MPORT_data = dataArray_7_9[dataArray_7_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_9_MPORT_addr = replace_set;
  assign dataArray_7_9_MPORT_mask = _GEN_1776 & _GEN_1571;
  assign dataArray_7_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_10_cachedata_MPORT_en = dataArray_7_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_10_cachedata_MPORT_addr = dataArray_7_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_10_cachedata_MPORT_data = dataArray_7_10[dataArray_7_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_10_MPORT_addr = replace_set;
  assign dataArray_7_10_MPORT_mask = _GEN_1776 & _GEN_1573;
  assign dataArray_7_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_11_cachedata_MPORT_en = dataArray_7_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_11_cachedata_MPORT_addr = dataArray_7_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_11_cachedata_MPORT_data = dataArray_7_11[dataArray_7_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_11_MPORT_addr = replace_set;
  assign dataArray_7_11_MPORT_mask = _GEN_1776 & _GEN_1575;
  assign dataArray_7_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_12_cachedata_MPORT_en = dataArray_7_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_12_cachedata_MPORT_addr = dataArray_7_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_12_cachedata_MPORT_data = dataArray_7_12[dataArray_7_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_12_MPORT_addr = replace_set;
  assign dataArray_7_12_MPORT_mask = _GEN_1776 & _GEN_1577;
  assign dataArray_7_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_13_cachedata_MPORT_en = dataArray_7_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_13_cachedata_MPORT_addr = dataArray_7_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_13_cachedata_MPORT_data = dataArray_7_13[dataArray_7_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_13_MPORT_addr = replace_set;
  assign dataArray_7_13_MPORT_mask = _GEN_1776 & _GEN_1579;
  assign dataArray_7_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_14_cachedata_MPORT_en = dataArray_7_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_14_cachedata_MPORT_addr = dataArray_7_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_14_cachedata_MPORT_data = dataArray_7_14[dataArray_7_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_14_MPORT_addr = replace_set;
  assign dataArray_7_14_MPORT_mask = _GEN_1776 & _GEN_1581;
  assign dataArray_7_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_7_15_cachedata_MPORT_en = dataArray_7_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_7_15_cachedata_MPORT_addr = dataArray_7_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_7_15_cachedata_MPORT_data = dataArray_7_15[dataArray_7_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_7_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_7_15_MPORT_addr = replace_set;
  assign dataArray_7_15_MPORT_mask = _GEN_1776 & _GEN_1583;
  assign dataArray_7_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_0_cachedata_MPORT_en = dataArray_8_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_0_cachedata_MPORT_addr = dataArray_8_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_0_cachedata_MPORT_data = dataArray_8_0[dataArray_8_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_0_MPORT_addr = replace_set;
  assign dataArray_8_0_MPORT_mask = _GEN_1808 & _GEN_1553;
  assign dataArray_8_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_1_cachedata_MPORT_en = dataArray_8_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_1_cachedata_MPORT_addr = dataArray_8_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_1_cachedata_MPORT_data = dataArray_8_1[dataArray_8_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_1_MPORT_addr = replace_set;
  assign dataArray_8_1_MPORT_mask = _GEN_1808 & _GEN_1555;
  assign dataArray_8_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_2_cachedata_MPORT_en = dataArray_8_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_2_cachedata_MPORT_addr = dataArray_8_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_2_cachedata_MPORT_data = dataArray_8_2[dataArray_8_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_2_MPORT_addr = replace_set;
  assign dataArray_8_2_MPORT_mask = _GEN_1808 & _GEN_1557;
  assign dataArray_8_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_3_cachedata_MPORT_en = dataArray_8_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_3_cachedata_MPORT_addr = dataArray_8_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_3_cachedata_MPORT_data = dataArray_8_3[dataArray_8_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_3_MPORT_addr = replace_set;
  assign dataArray_8_3_MPORT_mask = _GEN_1808 & _GEN_1559;
  assign dataArray_8_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_4_cachedata_MPORT_en = dataArray_8_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_4_cachedata_MPORT_addr = dataArray_8_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_4_cachedata_MPORT_data = dataArray_8_4[dataArray_8_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_4_MPORT_addr = replace_set;
  assign dataArray_8_4_MPORT_mask = _GEN_1808 & _GEN_1561;
  assign dataArray_8_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_5_cachedata_MPORT_en = dataArray_8_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_5_cachedata_MPORT_addr = dataArray_8_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_5_cachedata_MPORT_data = dataArray_8_5[dataArray_8_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_5_MPORT_addr = replace_set;
  assign dataArray_8_5_MPORT_mask = _GEN_1808 & _GEN_1563;
  assign dataArray_8_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_6_cachedata_MPORT_en = dataArray_8_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_6_cachedata_MPORT_addr = dataArray_8_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_6_cachedata_MPORT_data = dataArray_8_6[dataArray_8_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_6_MPORT_addr = replace_set;
  assign dataArray_8_6_MPORT_mask = _GEN_1808 & _GEN_1565;
  assign dataArray_8_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_7_cachedata_MPORT_en = dataArray_8_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_7_cachedata_MPORT_addr = dataArray_8_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_7_cachedata_MPORT_data = dataArray_8_7[dataArray_8_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_7_MPORT_addr = replace_set;
  assign dataArray_8_7_MPORT_mask = _GEN_1808 & _GEN_1567;
  assign dataArray_8_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_8_cachedata_MPORT_en = dataArray_8_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_8_cachedata_MPORT_addr = dataArray_8_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_8_cachedata_MPORT_data = dataArray_8_8[dataArray_8_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_8_MPORT_addr = replace_set;
  assign dataArray_8_8_MPORT_mask = _GEN_1808 & _GEN_1569;
  assign dataArray_8_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_9_cachedata_MPORT_en = dataArray_8_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_9_cachedata_MPORT_addr = dataArray_8_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_9_cachedata_MPORT_data = dataArray_8_9[dataArray_8_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_9_MPORT_addr = replace_set;
  assign dataArray_8_9_MPORT_mask = _GEN_1808 & _GEN_1571;
  assign dataArray_8_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_10_cachedata_MPORT_en = dataArray_8_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_10_cachedata_MPORT_addr = dataArray_8_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_10_cachedata_MPORT_data = dataArray_8_10[dataArray_8_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_10_MPORT_addr = replace_set;
  assign dataArray_8_10_MPORT_mask = _GEN_1808 & _GEN_1573;
  assign dataArray_8_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_11_cachedata_MPORT_en = dataArray_8_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_11_cachedata_MPORT_addr = dataArray_8_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_11_cachedata_MPORT_data = dataArray_8_11[dataArray_8_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_11_MPORT_addr = replace_set;
  assign dataArray_8_11_MPORT_mask = _GEN_1808 & _GEN_1575;
  assign dataArray_8_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_12_cachedata_MPORT_en = dataArray_8_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_12_cachedata_MPORT_addr = dataArray_8_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_12_cachedata_MPORT_data = dataArray_8_12[dataArray_8_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_12_MPORT_addr = replace_set;
  assign dataArray_8_12_MPORT_mask = _GEN_1808 & _GEN_1577;
  assign dataArray_8_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_13_cachedata_MPORT_en = dataArray_8_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_13_cachedata_MPORT_addr = dataArray_8_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_13_cachedata_MPORT_data = dataArray_8_13[dataArray_8_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_13_MPORT_addr = replace_set;
  assign dataArray_8_13_MPORT_mask = _GEN_1808 & _GEN_1579;
  assign dataArray_8_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_14_cachedata_MPORT_en = dataArray_8_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_14_cachedata_MPORT_addr = dataArray_8_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_14_cachedata_MPORT_data = dataArray_8_14[dataArray_8_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_14_MPORT_addr = replace_set;
  assign dataArray_8_14_MPORT_mask = _GEN_1808 & _GEN_1581;
  assign dataArray_8_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_8_15_cachedata_MPORT_en = dataArray_8_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_8_15_cachedata_MPORT_addr = dataArray_8_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_8_15_cachedata_MPORT_data = dataArray_8_15[dataArray_8_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_8_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_8_15_MPORT_addr = replace_set;
  assign dataArray_8_15_MPORT_mask = _GEN_1808 & _GEN_1583;
  assign dataArray_8_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_0_cachedata_MPORT_en = dataArray_9_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_0_cachedata_MPORT_addr = dataArray_9_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_0_cachedata_MPORT_data = dataArray_9_0[dataArray_9_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_0_MPORT_addr = replace_set;
  assign dataArray_9_0_MPORT_mask = _GEN_1840 & _GEN_1553;
  assign dataArray_9_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_1_cachedata_MPORT_en = dataArray_9_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_1_cachedata_MPORT_addr = dataArray_9_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_1_cachedata_MPORT_data = dataArray_9_1[dataArray_9_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_1_MPORT_addr = replace_set;
  assign dataArray_9_1_MPORT_mask = _GEN_1840 & _GEN_1555;
  assign dataArray_9_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_2_cachedata_MPORT_en = dataArray_9_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_2_cachedata_MPORT_addr = dataArray_9_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_2_cachedata_MPORT_data = dataArray_9_2[dataArray_9_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_2_MPORT_addr = replace_set;
  assign dataArray_9_2_MPORT_mask = _GEN_1840 & _GEN_1557;
  assign dataArray_9_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_3_cachedata_MPORT_en = dataArray_9_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_3_cachedata_MPORT_addr = dataArray_9_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_3_cachedata_MPORT_data = dataArray_9_3[dataArray_9_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_3_MPORT_addr = replace_set;
  assign dataArray_9_3_MPORT_mask = _GEN_1840 & _GEN_1559;
  assign dataArray_9_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_4_cachedata_MPORT_en = dataArray_9_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_4_cachedata_MPORT_addr = dataArray_9_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_4_cachedata_MPORT_data = dataArray_9_4[dataArray_9_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_4_MPORT_addr = replace_set;
  assign dataArray_9_4_MPORT_mask = _GEN_1840 & _GEN_1561;
  assign dataArray_9_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_5_cachedata_MPORT_en = dataArray_9_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_5_cachedata_MPORT_addr = dataArray_9_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_5_cachedata_MPORT_data = dataArray_9_5[dataArray_9_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_5_MPORT_addr = replace_set;
  assign dataArray_9_5_MPORT_mask = _GEN_1840 & _GEN_1563;
  assign dataArray_9_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_6_cachedata_MPORT_en = dataArray_9_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_6_cachedata_MPORT_addr = dataArray_9_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_6_cachedata_MPORT_data = dataArray_9_6[dataArray_9_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_6_MPORT_addr = replace_set;
  assign dataArray_9_6_MPORT_mask = _GEN_1840 & _GEN_1565;
  assign dataArray_9_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_7_cachedata_MPORT_en = dataArray_9_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_7_cachedata_MPORT_addr = dataArray_9_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_7_cachedata_MPORT_data = dataArray_9_7[dataArray_9_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_7_MPORT_addr = replace_set;
  assign dataArray_9_7_MPORT_mask = _GEN_1840 & _GEN_1567;
  assign dataArray_9_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_8_cachedata_MPORT_en = dataArray_9_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_8_cachedata_MPORT_addr = dataArray_9_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_8_cachedata_MPORT_data = dataArray_9_8[dataArray_9_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_8_MPORT_addr = replace_set;
  assign dataArray_9_8_MPORT_mask = _GEN_1840 & _GEN_1569;
  assign dataArray_9_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_9_cachedata_MPORT_en = dataArray_9_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_9_cachedata_MPORT_addr = dataArray_9_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_9_cachedata_MPORT_data = dataArray_9_9[dataArray_9_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_9_MPORT_addr = replace_set;
  assign dataArray_9_9_MPORT_mask = _GEN_1840 & _GEN_1571;
  assign dataArray_9_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_10_cachedata_MPORT_en = dataArray_9_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_10_cachedata_MPORT_addr = dataArray_9_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_10_cachedata_MPORT_data = dataArray_9_10[dataArray_9_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_10_MPORT_addr = replace_set;
  assign dataArray_9_10_MPORT_mask = _GEN_1840 & _GEN_1573;
  assign dataArray_9_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_11_cachedata_MPORT_en = dataArray_9_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_11_cachedata_MPORT_addr = dataArray_9_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_11_cachedata_MPORT_data = dataArray_9_11[dataArray_9_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_11_MPORT_addr = replace_set;
  assign dataArray_9_11_MPORT_mask = _GEN_1840 & _GEN_1575;
  assign dataArray_9_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_12_cachedata_MPORT_en = dataArray_9_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_12_cachedata_MPORT_addr = dataArray_9_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_12_cachedata_MPORT_data = dataArray_9_12[dataArray_9_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_12_MPORT_addr = replace_set;
  assign dataArray_9_12_MPORT_mask = _GEN_1840 & _GEN_1577;
  assign dataArray_9_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_13_cachedata_MPORT_en = dataArray_9_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_13_cachedata_MPORT_addr = dataArray_9_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_13_cachedata_MPORT_data = dataArray_9_13[dataArray_9_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_13_MPORT_addr = replace_set;
  assign dataArray_9_13_MPORT_mask = _GEN_1840 & _GEN_1579;
  assign dataArray_9_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_14_cachedata_MPORT_en = dataArray_9_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_14_cachedata_MPORT_addr = dataArray_9_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_14_cachedata_MPORT_data = dataArray_9_14[dataArray_9_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_14_MPORT_addr = replace_set;
  assign dataArray_9_14_MPORT_mask = _GEN_1840 & _GEN_1581;
  assign dataArray_9_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_9_15_cachedata_MPORT_en = dataArray_9_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_9_15_cachedata_MPORT_addr = dataArray_9_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_9_15_cachedata_MPORT_data = dataArray_9_15[dataArray_9_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_9_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_9_15_MPORT_addr = replace_set;
  assign dataArray_9_15_MPORT_mask = _GEN_1840 & _GEN_1583;
  assign dataArray_9_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_0_cachedata_MPORT_en = dataArray_10_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_0_cachedata_MPORT_addr = dataArray_10_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_0_cachedata_MPORT_data = dataArray_10_0[dataArray_10_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_0_MPORT_addr = replace_set;
  assign dataArray_10_0_MPORT_mask = _GEN_1872 & _GEN_1553;
  assign dataArray_10_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_1_cachedata_MPORT_en = dataArray_10_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_1_cachedata_MPORT_addr = dataArray_10_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_1_cachedata_MPORT_data = dataArray_10_1[dataArray_10_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_1_MPORT_addr = replace_set;
  assign dataArray_10_1_MPORT_mask = _GEN_1872 & _GEN_1555;
  assign dataArray_10_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_2_cachedata_MPORT_en = dataArray_10_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_2_cachedata_MPORT_addr = dataArray_10_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_2_cachedata_MPORT_data = dataArray_10_2[dataArray_10_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_2_MPORT_addr = replace_set;
  assign dataArray_10_2_MPORT_mask = _GEN_1872 & _GEN_1557;
  assign dataArray_10_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_3_cachedata_MPORT_en = dataArray_10_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_3_cachedata_MPORT_addr = dataArray_10_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_3_cachedata_MPORT_data = dataArray_10_3[dataArray_10_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_3_MPORT_addr = replace_set;
  assign dataArray_10_3_MPORT_mask = _GEN_1872 & _GEN_1559;
  assign dataArray_10_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_4_cachedata_MPORT_en = dataArray_10_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_4_cachedata_MPORT_addr = dataArray_10_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_4_cachedata_MPORT_data = dataArray_10_4[dataArray_10_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_4_MPORT_addr = replace_set;
  assign dataArray_10_4_MPORT_mask = _GEN_1872 & _GEN_1561;
  assign dataArray_10_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_5_cachedata_MPORT_en = dataArray_10_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_5_cachedata_MPORT_addr = dataArray_10_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_5_cachedata_MPORT_data = dataArray_10_5[dataArray_10_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_5_MPORT_addr = replace_set;
  assign dataArray_10_5_MPORT_mask = _GEN_1872 & _GEN_1563;
  assign dataArray_10_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_6_cachedata_MPORT_en = dataArray_10_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_6_cachedata_MPORT_addr = dataArray_10_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_6_cachedata_MPORT_data = dataArray_10_6[dataArray_10_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_6_MPORT_addr = replace_set;
  assign dataArray_10_6_MPORT_mask = _GEN_1872 & _GEN_1565;
  assign dataArray_10_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_7_cachedata_MPORT_en = dataArray_10_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_7_cachedata_MPORT_addr = dataArray_10_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_7_cachedata_MPORT_data = dataArray_10_7[dataArray_10_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_7_MPORT_addr = replace_set;
  assign dataArray_10_7_MPORT_mask = _GEN_1872 & _GEN_1567;
  assign dataArray_10_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_8_cachedata_MPORT_en = dataArray_10_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_8_cachedata_MPORT_addr = dataArray_10_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_8_cachedata_MPORT_data = dataArray_10_8[dataArray_10_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_8_MPORT_addr = replace_set;
  assign dataArray_10_8_MPORT_mask = _GEN_1872 & _GEN_1569;
  assign dataArray_10_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_9_cachedata_MPORT_en = dataArray_10_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_9_cachedata_MPORT_addr = dataArray_10_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_9_cachedata_MPORT_data = dataArray_10_9[dataArray_10_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_9_MPORT_addr = replace_set;
  assign dataArray_10_9_MPORT_mask = _GEN_1872 & _GEN_1571;
  assign dataArray_10_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_10_cachedata_MPORT_en = dataArray_10_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_10_cachedata_MPORT_addr = dataArray_10_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_10_cachedata_MPORT_data = dataArray_10_10[dataArray_10_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_10_MPORT_addr = replace_set;
  assign dataArray_10_10_MPORT_mask = _GEN_1872 & _GEN_1573;
  assign dataArray_10_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_11_cachedata_MPORT_en = dataArray_10_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_11_cachedata_MPORT_addr = dataArray_10_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_11_cachedata_MPORT_data = dataArray_10_11[dataArray_10_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_11_MPORT_addr = replace_set;
  assign dataArray_10_11_MPORT_mask = _GEN_1872 & _GEN_1575;
  assign dataArray_10_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_12_cachedata_MPORT_en = dataArray_10_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_12_cachedata_MPORT_addr = dataArray_10_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_12_cachedata_MPORT_data = dataArray_10_12[dataArray_10_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_12_MPORT_addr = replace_set;
  assign dataArray_10_12_MPORT_mask = _GEN_1872 & _GEN_1577;
  assign dataArray_10_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_13_cachedata_MPORT_en = dataArray_10_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_13_cachedata_MPORT_addr = dataArray_10_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_13_cachedata_MPORT_data = dataArray_10_13[dataArray_10_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_13_MPORT_addr = replace_set;
  assign dataArray_10_13_MPORT_mask = _GEN_1872 & _GEN_1579;
  assign dataArray_10_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_14_cachedata_MPORT_en = dataArray_10_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_14_cachedata_MPORT_addr = dataArray_10_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_14_cachedata_MPORT_data = dataArray_10_14[dataArray_10_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_14_MPORT_addr = replace_set;
  assign dataArray_10_14_MPORT_mask = _GEN_1872 & _GEN_1581;
  assign dataArray_10_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_10_15_cachedata_MPORT_en = dataArray_10_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_10_15_cachedata_MPORT_addr = dataArray_10_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_10_15_cachedata_MPORT_data = dataArray_10_15[dataArray_10_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_10_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_10_15_MPORT_addr = replace_set;
  assign dataArray_10_15_MPORT_mask = _GEN_1872 & _GEN_1583;
  assign dataArray_10_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_0_cachedata_MPORT_en = dataArray_11_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_0_cachedata_MPORT_addr = dataArray_11_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_0_cachedata_MPORT_data = dataArray_11_0[dataArray_11_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_0_MPORT_addr = replace_set;
  assign dataArray_11_0_MPORT_mask = _GEN_1904 & _GEN_1553;
  assign dataArray_11_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_1_cachedata_MPORT_en = dataArray_11_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_1_cachedata_MPORT_addr = dataArray_11_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_1_cachedata_MPORT_data = dataArray_11_1[dataArray_11_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_1_MPORT_addr = replace_set;
  assign dataArray_11_1_MPORT_mask = _GEN_1904 & _GEN_1555;
  assign dataArray_11_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_2_cachedata_MPORT_en = dataArray_11_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_2_cachedata_MPORT_addr = dataArray_11_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_2_cachedata_MPORT_data = dataArray_11_2[dataArray_11_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_2_MPORT_addr = replace_set;
  assign dataArray_11_2_MPORT_mask = _GEN_1904 & _GEN_1557;
  assign dataArray_11_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_3_cachedata_MPORT_en = dataArray_11_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_3_cachedata_MPORT_addr = dataArray_11_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_3_cachedata_MPORT_data = dataArray_11_3[dataArray_11_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_3_MPORT_addr = replace_set;
  assign dataArray_11_3_MPORT_mask = _GEN_1904 & _GEN_1559;
  assign dataArray_11_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_4_cachedata_MPORT_en = dataArray_11_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_4_cachedata_MPORT_addr = dataArray_11_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_4_cachedata_MPORT_data = dataArray_11_4[dataArray_11_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_4_MPORT_addr = replace_set;
  assign dataArray_11_4_MPORT_mask = _GEN_1904 & _GEN_1561;
  assign dataArray_11_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_5_cachedata_MPORT_en = dataArray_11_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_5_cachedata_MPORT_addr = dataArray_11_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_5_cachedata_MPORT_data = dataArray_11_5[dataArray_11_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_5_MPORT_addr = replace_set;
  assign dataArray_11_5_MPORT_mask = _GEN_1904 & _GEN_1563;
  assign dataArray_11_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_6_cachedata_MPORT_en = dataArray_11_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_6_cachedata_MPORT_addr = dataArray_11_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_6_cachedata_MPORT_data = dataArray_11_6[dataArray_11_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_6_MPORT_addr = replace_set;
  assign dataArray_11_6_MPORT_mask = _GEN_1904 & _GEN_1565;
  assign dataArray_11_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_7_cachedata_MPORT_en = dataArray_11_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_7_cachedata_MPORT_addr = dataArray_11_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_7_cachedata_MPORT_data = dataArray_11_7[dataArray_11_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_7_MPORT_addr = replace_set;
  assign dataArray_11_7_MPORT_mask = _GEN_1904 & _GEN_1567;
  assign dataArray_11_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_8_cachedata_MPORT_en = dataArray_11_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_8_cachedata_MPORT_addr = dataArray_11_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_8_cachedata_MPORT_data = dataArray_11_8[dataArray_11_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_8_MPORT_addr = replace_set;
  assign dataArray_11_8_MPORT_mask = _GEN_1904 & _GEN_1569;
  assign dataArray_11_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_9_cachedata_MPORT_en = dataArray_11_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_9_cachedata_MPORT_addr = dataArray_11_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_9_cachedata_MPORT_data = dataArray_11_9[dataArray_11_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_9_MPORT_addr = replace_set;
  assign dataArray_11_9_MPORT_mask = _GEN_1904 & _GEN_1571;
  assign dataArray_11_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_10_cachedata_MPORT_en = dataArray_11_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_10_cachedata_MPORT_addr = dataArray_11_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_10_cachedata_MPORT_data = dataArray_11_10[dataArray_11_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_10_MPORT_addr = replace_set;
  assign dataArray_11_10_MPORT_mask = _GEN_1904 & _GEN_1573;
  assign dataArray_11_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_11_cachedata_MPORT_en = dataArray_11_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_11_cachedata_MPORT_addr = dataArray_11_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_11_cachedata_MPORT_data = dataArray_11_11[dataArray_11_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_11_MPORT_addr = replace_set;
  assign dataArray_11_11_MPORT_mask = _GEN_1904 & _GEN_1575;
  assign dataArray_11_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_12_cachedata_MPORT_en = dataArray_11_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_12_cachedata_MPORT_addr = dataArray_11_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_12_cachedata_MPORT_data = dataArray_11_12[dataArray_11_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_12_MPORT_addr = replace_set;
  assign dataArray_11_12_MPORT_mask = _GEN_1904 & _GEN_1577;
  assign dataArray_11_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_13_cachedata_MPORT_en = dataArray_11_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_13_cachedata_MPORT_addr = dataArray_11_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_13_cachedata_MPORT_data = dataArray_11_13[dataArray_11_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_13_MPORT_addr = replace_set;
  assign dataArray_11_13_MPORT_mask = _GEN_1904 & _GEN_1579;
  assign dataArray_11_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_14_cachedata_MPORT_en = dataArray_11_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_14_cachedata_MPORT_addr = dataArray_11_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_14_cachedata_MPORT_data = dataArray_11_14[dataArray_11_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_14_MPORT_addr = replace_set;
  assign dataArray_11_14_MPORT_mask = _GEN_1904 & _GEN_1581;
  assign dataArray_11_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_11_15_cachedata_MPORT_en = dataArray_11_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_11_15_cachedata_MPORT_addr = dataArray_11_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_11_15_cachedata_MPORT_data = dataArray_11_15[dataArray_11_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_11_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_11_15_MPORT_addr = replace_set;
  assign dataArray_11_15_MPORT_mask = _GEN_1904 & _GEN_1583;
  assign dataArray_11_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_0_cachedata_MPORT_en = dataArray_12_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_0_cachedata_MPORT_addr = dataArray_12_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_0_cachedata_MPORT_data = dataArray_12_0[dataArray_12_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_0_MPORT_addr = replace_set;
  assign dataArray_12_0_MPORT_mask = _GEN_1936 & _GEN_1553;
  assign dataArray_12_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_1_cachedata_MPORT_en = dataArray_12_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_1_cachedata_MPORT_addr = dataArray_12_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_1_cachedata_MPORT_data = dataArray_12_1[dataArray_12_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_1_MPORT_addr = replace_set;
  assign dataArray_12_1_MPORT_mask = _GEN_1936 & _GEN_1555;
  assign dataArray_12_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_2_cachedata_MPORT_en = dataArray_12_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_2_cachedata_MPORT_addr = dataArray_12_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_2_cachedata_MPORT_data = dataArray_12_2[dataArray_12_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_2_MPORT_addr = replace_set;
  assign dataArray_12_2_MPORT_mask = _GEN_1936 & _GEN_1557;
  assign dataArray_12_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_3_cachedata_MPORT_en = dataArray_12_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_3_cachedata_MPORT_addr = dataArray_12_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_3_cachedata_MPORT_data = dataArray_12_3[dataArray_12_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_3_MPORT_addr = replace_set;
  assign dataArray_12_3_MPORT_mask = _GEN_1936 & _GEN_1559;
  assign dataArray_12_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_4_cachedata_MPORT_en = dataArray_12_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_4_cachedata_MPORT_addr = dataArray_12_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_4_cachedata_MPORT_data = dataArray_12_4[dataArray_12_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_4_MPORT_addr = replace_set;
  assign dataArray_12_4_MPORT_mask = _GEN_1936 & _GEN_1561;
  assign dataArray_12_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_5_cachedata_MPORT_en = dataArray_12_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_5_cachedata_MPORT_addr = dataArray_12_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_5_cachedata_MPORT_data = dataArray_12_5[dataArray_12_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_5_MPORT_addr = replace_set;
  assign dataArray_12_5_MPORT_mask = _GEN_1936 & _GEN_1563;
  assign dataArray_12_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_6_cachedata_MPORT_en = dataArray_12_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_6_cachedata_MPORT_addr = dataArray_12_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_6_cachedata_MPORT_data = dataArray_12_6[dataArray_12_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_6_MPORT_addr = replace_set;
  assign dataArray_12_6_MPORT_mask = _GEN_1936 & _GEN_1565;
  assign dataArray_12_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_7_cachedata_MPORT_en = dataArray_12_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_7_cachedata_MPORT_addr = dataArray_12_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_7_cachedata_MPORT_data = dataArray_12_7[dataArray_12_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_7_MPORT_addr = replace_set;
  assign dataArray_12_7_MPORT_mask = _GEN_1936 & _GEN_1567;
  assign dataArray_12_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_8_cachedata_MPORT_en = dataArray_12_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_8_cachedata_MPORT_addr = dataArray_12_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_8_cachedata_MPORT_data = dataArray_12_8[dataArray_12_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_8_MPORT_addr = replace_set;
  assign dataArray_12_8_MPORT_mask = _GEN_1936 & _GEN_1569;
  assign dataArray_12_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_9_cachedata_MPORT_en = dataArray_12_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_9_cachedata_MPORT_addr = dataArray_12_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_9_cachedata_MPORT_data = dataArray_12_9[dataArray_12_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_9_MPORT_addr = replace_set;
  assign dataArray_12_9_MPORT_mask = _GEN_1936 & _GEN_1571;
  assign dataArray_12_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_10_cachedata_MPORT_en = dataArray_12_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_10_cachedata_MPORT_addr = dataArray_12_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_10_cachedata_MPORT_data = dataArray_12_10[dataArray_12_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_10_MPORT_addr = replace_set;
  assign dataArray_12_10_MPORT_mask = _GEN_1936 & _GEN_1573;
  assign dataArray_12_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_11_cachedata_MPORT_en = dataArray_12_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_11_cachedata_MPORT_addr = dataArray_12_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_11_cachedata_MPORT_data = dataArray_12_11[dataArray_12_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_11_MPORT_addr = replace_set;
  assign dataArray_12_11_MPORT_mask = _GEN_1936 & _GEN_1575;
  assign dataArray_12_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_12_cachedata_MPORT_en = dataArray_12_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_12_cachedata_MPORT_addr = dataArray_12_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_12_cachedata_MPORT_data = dataArray_12_12[dataArray_12_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_12_MPORT_addr = replace_set;
  assign dataArray_12_12_MPORT_mask = _GEN_1936 & _GEN_1577;
  assign dataArray_12_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_13_cachedata_MPORT_en = dataArray_12_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_13_cachedata_MPORT_addr = dataArray_12_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_13_cachedata_MPORT_data = dataArray_12_13[dataArray_12_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_13_MPORT_addr = replace_set;
  assign dataArray_12_13_MPORT_mask = _GEN_1936 & _GEN_1579;
  assign dataArray_12_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_14_cachedata_MPORT_en = dataArray_12_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_14_cachedata_MPORT_addr = dataArray_12_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_14_cachedata_MPORT_data = dataArray_12_14[dataArray_12_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_14_MPORT_addr = replace_set;
  assign dataArray_12_14_MPORT_mask = _GEN_1936 & _GEN_1581;
  assign dataArray_12_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_12_15_cachedata_MPORT_en = dataArray_12_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_12_15_cachedata_MPORT_addr = dataArray_12_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_12_15_cachedata_MPORT_data = dataArray_12_15[dataArray_12_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_12_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_12_15_MPORT_addr = replace_set;
  assign dataArray_12_15_MPORT_mask = _GEN_1936 & _GEN_1583;
  assign dataArray_12_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_0_cachedata_MPORT_en = dataArray_13_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_0_cachedata_MPORT_addr = dataArray_13_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_0_cachedata_MPORT_data = dataArray_13_0[dataArray_13_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_0_MPORT_addr = replace_set;
  assign dataArray_13_0_MPORT_mask = _GEN_1968 & _GEN_1553;
  assign dataArray_13_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_1_cachedata_MPORT_en = dataArray_13_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_1_cachedata_MPORT_addr = dataArray_13_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_1_cachedata_MPORT_data = dataArray_13_1[dataArray_13_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_1_MPORT_addr = replace_set;
  assign dataArray_13_1_MPORT_mask = _GEN_1968 & _GEN_1555;
  assign dataArray_13_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_2_cachedata_MPORT_en = dataArray_13_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_2_cachedata_MPORT_addr = dataArray_13_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_2_cachedata_MPORT_data = dataArray_13_2[dataArray_13_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_2_MPORT_addr = replace_set;
  assign dataArray_13_2_MPORT_mask = _GEN_1968 & _GEN_1557;
  assign dataArray_13_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_3_cachedata_MPORT_en = dataArray_13_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_3_cachedata_MPORT_addr = dataArray_13_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_3_cachedata_MPORT_data = dataArray_13_3[dataArray_13_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_3_MPORT_addr = replace_set;
  assign dataArray_13_3_MPORT_mask = _GEN_1968 & _GEN_1559;
  assign dataArray_13_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_4_cachedata_MPORT_en = dataArray_13_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_4_cachedata_MPORT_addr = dataArray_13_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_4_cachedata_MPORT_data = dataArray_13_4[dataArray_13_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_4_MPORT_addr = replace_set;
  assign dataArray_13_4_MPORT_mask = _GEN_1968 & _GEN_1561;
  assign dataArray_13_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_5_cachedata_MPORT_en = dataArray_13_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_5_cachedata_MPORT_addr = dataArray_13_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_5_cachedata_MPORT_data = dataArray_13_5[dataArray_13_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_5_MPORT_addr = replace_set;
  assign dataArray_13_5_MPORT_mask = _GEN_1968 & _GEN_1563;
  assign dataArray_13_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_6_cachedata_MPORT_en = dataArray_13_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_6_cachedata_MPORT_addr = dataArray_13_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_6_cachedata_MPORT_data = dataArray_13_6[dataArray_13_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_6_MPORT_addr = replace_set;
  assign dataArray_13_6_MPORT_mask = _GEN_1968 & _GEN_1565;
  assign dataArray_13_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_7_cachedata_MPORT_en = dataArray_13_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_7_cachedata_MPORT_addr = dataArray_13_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_7_cachedata_MPORT_data = dataArray_13_7[dataArray_13_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_7_MPORT_addr = replace_set;
  assign dataArray_13_7_MPORT_mask = _GEN_1968 & _GEN_1567;
  assign dataArray_13_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_8_cachedata_MPORT_en = dataArray_13_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_8_cachedata_MPORT_addr = dataArray_13_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_8_cachedata_MPORT_data = dataArray_13_8[dataArray_13_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_8_MPORT_addr = replace_set;
  assign dataArray_13_8_MPORT_mask = _GEN_1968 & _GEN_1569;
  assign dataArray_13_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_9_cachedata_MPORT_en = dataArray_13_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_9_cachedata_MPORT_addr = dataArray_13_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_9_cachedata_MPORT_data = dataArray_13_9[dataArray_13_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_9_MPORT_addr = replace_set;
  assign dataArray_13_9_MPORT_mask = _GEN_1968 & _GEN_1571;
  assign dataArray_13_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_10_cachedata_MPORT_en = dataArray_13_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_10_cachedata_MPORT_addr = dataArray_13_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_10_cachedata_MPORT_data = dataArray_13_10[dataArray_13_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_10_MPORT_addr = replace_set;
  assign dataArray_13_10_MPORT_mask = _GEN_1968 & _GEN_1573;
  assign dataArray_13_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_11_cachedata_MPORT_en = dataArray_13_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_11_cachedata_MPORT_addr = dataArray_13_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_11_cachedata_MPORT_data = dataArray_13_11[dataArray_13_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_11_MPORT_addr = replace_set;
  assign dataArray_13_11_MPORT_mask = _GEN_1968 & _GEN_1575;
  assign dataArray_13_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_12_cachedata_MPORT_en = dataArray_13_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_12_cachedata_MPORT_addr = dataArray_13_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_12_cachedata_MPORT_data = dataArray_13_12[dataArray_13_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_12_MPORT_addr = replace_set;
  assign dataArray_13_12_MPORT_mask = _GEN_1968 & _GEN_1577;
  assign dataArray_13_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_13_cachedata_MPORT_en = dataArray_13_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_13_cachedata_MPORT_addr = dataArray_13_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_13_cachedata_MPORT_data = dataArray_13_13[dataArray_13_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_13_MPORT_addr = replace_set;
  assign dataArray_13_13_MPORT_mask = _GEN_1968 & _GEN_1579;
  assign dataArray_13_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_14_cachedata_MPORT_en = dataArray_13_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_14_cachedata_MPORT_addr = dataArray_13_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_14_cachedata_MPORT_data = dataArray_13_14[dataArray_13_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_14_MPORT_addr = replace_set;
  assign dataArray_13_14_MPORT_mask = _GEN_1968 & _GEN_1581;
  assign dataArray_13_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_13_15_cachedata_MPORT_en = dataArray_13_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_13_15_cachedata_MPORT_addr = dataArray_13_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_13_15_cachedata_MPORT_data = dataArray_13_15[dataArray_13_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_13_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_13_15_MPORT_addr = replace_set;
  assign dataArray_13_15_MPORT_mask = _GEN_1968 & _GEN_1583;
  assign dataArray_13_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_0_cachedata_MPORT_en = dataArray_14_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_0_cachedata_MPORT_addr = dataArray_14_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_0_cachedata_MPORT_data = dataArray_14_0[dataArray_14_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_0_MPORT_addr = replace_set;
  assign dataArray_14_0_MPORT_mask = _GEN_2000 & _GEN_1553;
  assign dataArray_14_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_1_cachedata_MPORT_en = dataArray_14_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_1_cachedata_MPORT_addr = dataArray_14_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_1_cachedata_MPORT_data = dataArray_14_1[dataArray_14_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_1_MPORT_addr = replace_set;
  assign dataArray_14_1_MPORT_mask = _GEN_2000 & _GEN_1555;
  assign dataArray_14_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_2_cachedata_MPORT_en = dataArray_14_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_2_cachedata_MPORT_addr = dataArray_14_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_2_cachedata_MPORT_data = dataArray_14_2[dataArray_14_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_2_MPORT_addr = replace_set;
  assign dataArray_14_2_MPORT_mask = _GEN_2000 & _GEN_1557;
  assign dataArray_14_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_3_cachedata_MPORT_en = dataArray_14_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_3_cachedata_MPORT_addr = dataArray_14_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_3_cachedata_MPORT_data = dataArray_14_3[dataArray_14_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_3_MPORT_addr = replace_set;
  assign dataArray_14_3_MPORT_mask = _GEN_2000 & _GEN_1559;
  assign dataArray_14_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_4_cachedata_MPORT_en = dataArray_14_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_4_cachedata_MPORT_addr = dataArray_14_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_4_cachedata_MPORT_data = dataArray_14_4[dataArray_14_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_4_MPORT_addr = replace_set;
  assign dataArray_14_4_MPORT_mask = _GEN_2000 & _GEN_1561;
  assign dataArray_14_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_5_cachedata_MPORT_en = dataArray_14_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_5_cachedata_MPORT_addr = dataArray_14_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_5_cachedata_MPORT_data = dataArray_14_5[dataArray_14_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_5_MPORT_addr = replace_set;
  assign dataArray_14_5_MPORT_mask = _GEN_2000 & _GEN_1563;
  assign dataArray_14_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_6_cachedata_MPORT_en = dataArray_14_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_6_cachedata_MPORT_addr = dataArray_14_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_6_cachedata_MPORT_data = dataArray_14_6[dataArray_14_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_6_MPORT_addr = replace_set;
  assign dataArray_14_6_MPORT_mask = _GEN_2000 & _GEN_1565;
  assign dataArray_14_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_7_cachedata_MPORT_en = dataArray_14_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_7_cachedata_MPORT_addr = dataArray_14_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_7_cachedata_MPORT_data = dataArray_14_7[dataArray_14_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_7_MPORT_addr = replace_set;
  assign dataArray_14_7_MPORT_mask = _GEN_2000 & _GEN_1567;
  assign dataArray_14_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_8_cachedata_MPORT_en = dataArray_14_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_8_cachedata_MPORT_addr = dataArray_14_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_8_cachedata_MPORT_data = dataArray_14_8[dataArray_14_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_8_MPORT_addr = replace_set;
  assign dataArray_14_8_MPORT_mask = _GEN_2000 & _GEN_1569;
  assign dataArray_14_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_9_cachedata_MPORT_en = dataArray_14_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_9_cachedata_MPORT_addr = dataArray_14_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_9_cachedata_MPORT_data = dataArray_14_9[dataArray_14_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_9_MPORT_addr = replace_set;
  assign dataArray_14_9_MPORT_mask = _GEN_2000 & _GEN_1571;
  assign dataArray_14_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_10_cachedata_MPORT_en = dataArray_14_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_10_cachedata_MPORT_addr = dataArray_14_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_10_cachedata_MPORT_data = dataArray_14_10[dataArray_14_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_10_MPORT_addr = replace_set;
  assign dataArray_14_10_MPORT_mask = _GEN_2000 & _GEN_1573;
  assign dataArray_14_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_11_cachedata_MPORT_en = dataArray_14_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_11_cachedata_MPORT_addr = dataArray_14_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_11_cachedata_MPORT_data = dataArray_14_11[dataArray_14_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_11_MPORT_addr = replace_set;
  assign dataArray_14_11_MPORT_mask = _GEN_2000 & _GEN_1575;
  assign dataArray_14_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_12_cachedata_MPORT_en = dataArray_14_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_12_cachedata_MPORT_addr = dataArray_14_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_12_cachedata_MPORT_data = dataArray_14_12[dataArray_14_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_12_MPORT_addr = replace_set;
  assign dataArray_14_12_MPORT_mask = _GEN_2000 & _GEN_1577;
  assign dataArray_14_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_13_cachedata_MPORT_en = dataArray_14_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_13_cachedata_MPORT_addr = dataArray_14_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_13_cachedata_MPORT_data = dataArray_14_13[dataArray_14_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_13_MPORT_addr = replace_set;
  assign dataArray_14_13_MPORT_mask = _GEN_2000 & _GEN_1579;
  assign dataArray_14_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_14_cachedata_MPORT_en = dataArray_14_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_14_cachedata_MPORT_addr = dataArray_14_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_14_cachedata_MPORT_data = dataArray_14_14[dataArray_14_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_14_MPORT_addr = replace_set;
  assign dataArray_14_14_MPORT_mask = _GEN_2000 & _GEN_1581;
  assign dataArray_14_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_14_15_cachedata_MPORT_en = dataArray_14_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_14_15_cachedata_MPORT_addr = dataArray_14_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_14_15_cachedata_MPORT_data = dataArray_14_15[dataArray_14_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_14_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_14_15_MPORT_addr = replace_set;
  assign dataArray_14_15_MPORT_mask = _GEN_2000 & _GEN_1583;
  assign dataArray_14_15_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_0_cachedata_MPORT_en = dataArray_15_0_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_0_cachedata_MPORT_addr = dataArray_15_0_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_0_cachedata_MPORT_data = dataArray_15_0[dataArray_15_0_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_0_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_0_MPORT_addr = replace_set;
  assign dataArray_15_0_MPORT_mask = _GEN_2032 & _GEN_1553;
  assign dataArray_15_0_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_1_cachedata_MPORT_en = dataArray_15_1_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_1_cachedata_MPORT_addr = dataArray_15_1_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_1_cachedata_MPORT_data = dataArray_15_1[dataArray_15_1_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_1_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_1_MPORT_addr = replace_set;
  assign dataArray_15_1_MPORT_mask = _GEN_2032 & _GEN_1555;
  assign dataArray_15_1_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_2_cachedata_MPORT_en = dataArray_15_2_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_2_cachedata_MPORT_addr = dataArray_15_2_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_2_cachedata_MPORT_data = dataArray_15_2[dataArray_15_2_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_2_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_2_MPORT_addr = replace_set;
  assign dataArray_15_2_MPORT_mask = _GEN_2032 & _GEN_1557;
  assign dataArray_15_2_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_3_cachedata_MPORT_en = dataArray_15_3_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_3_cachedata_MPORT_addr = dataArray_15_3_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_3_cachedata_MPORT_data = dataArray_15_3[dataArray_15_3_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_3_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_3_MPORT_addr = replace_set;
  assign dataArray_15_3_MPORT_mask = _GEN_2032 & _GEN_1559;
  assign dataArray_15_3_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_4_cachedata_MPORT_en = dataArray_15_4_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_4_cachedata_MPORT_addr = dataArray_15_4_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_4_cachedata_MPORT_data = dataArray_15_4[dataArray_15_4_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_4_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_4_MPORT_addr = replace_set;
  assign dataArray_15_4_MPORT_mask = _GEN_2032 & _GEN_1561;
  assign dataArray_15_4_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_5_cachedata_MPORT_en = dataArray_15_5_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_5_cachedata_MPORT_addr = dataArray_15_5_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_5_cachedata_MPORT_data = dataArray_15_5[dataArray_15_5_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_5_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_5_MPORT_addr = replace_set;
  assign dataArray_15_5_MPORT_mask = _GEN_2032 & _GEN_1563;
  assign dataArray_15_5_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_6_cachedata_MPORT_en = dataArray_15_6_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_6_cachedata_MPORT_addr = dataArray_15_6_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_6_cachedata_MPORT_data = dataArray_15_6[dataArray_15_6_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_6_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_6_MPORT_addr = replace_set;
  assign dataArray_15_6_MPORT_mask = _GEN_2032 & _GEN_1565;
  assign dataArray_15_6_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_7_cachedata_MPORT_en = dataArray_15_7_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_7_cachedata_MPORT_addr = dataArray_15_7_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_7_cachedata_MPORT_data = dataArray_15_7[dataArray_15_7_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_7_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_7_MPORT_addr = replace_set;
  assign dataArray_15_7_MPORT_mask = _GEN_2032 & _GEN_1567;
  assign dataArray_15_7_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_8_cachedata_MPORT_en = dataArray_15_8_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_8_cachedata_MPORT_addr = dataArray_15_8_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_8_cachedata_MPORT_data = dataArray_15_8[dataArray_15_8_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_8_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_8_MPORT_addr = replace_set;
  assign dataArray_15_8_MPORT_mask = _GEN_2032 & _GEN_1569;
  assign dataArray_15_8_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_9_cachedata_MPORT_en = dataArray_15_9_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_9_cachedata_MPORT_addr = dataArray_15_9_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_9_cachedata_MPORT_data = dataArray_15_9[dataArray_15_9_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_9_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_9_MPORT_addr = replace_set;
  assign dataArray_15_9_MPORT_mask = _GEN_2032 & _GEN_1571;
  assign dataArray_15_9_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_10_cachedata_MPORT_en = dataArray_15_10_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_10_cachedata_MPORT_addr = dataArray_15_10_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_10_cachedata_MPORT_data = dataArray_15_10[dataArray_15_10_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_10_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_10_MPORT_addr = replace_set;
  assign dataArray_15_10_MPORT_mask = _GEN_2032 & _GEN_1573;
  assign dataArray_15_10_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_11_cachedata_MPORT_en = dataArray_15_11_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_11_cachedata_MPORT_addr = dataArray_15_11_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_11_cachedata_MPORT_data = dataArray_15_11[dataArray_15_11_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_11_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_11_MPORT_addr = replace_set;
  assign dataArray_15_11_MPORT_mask = _GEN_2032 & _GEN_1575;
  assign dataArray_15_11_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_12_cachedata_MPORT_en = dataArray_15_12_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_12_cachedata_MPORT_addr = dataArray_15_12_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_12_cachedata_MPORT_data = dataArray_15_12[dataArray_15_12_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_12_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_12_MPORT_addr = replace_set;
  assign dataArray_15_12_MPORT_mask = _GEN_2032 & _GEN_1577;
  assign dataArray_15_12_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_13_cachedata_MPORT_en = dataArray_15_13_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_13_cachedata_MPORT_addr = dataArray_15_13_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_13_cachedata_MPORT_data = dataArray_15_13[dataArray_15_13_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_13_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_13_MPORT_addr = replace_set;
  assign dataArray_15_13_MPORT_mask = _GEN_2032 & _GEN_1579;
  assign dataArray_15_13_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_14_cachedata_MPORT_en = dataArray_15_14_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_14_cachedata_MPORT_addr = dataArray_15_14_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_14_cachedata_MPORT_data = dataArray_15_14[dataArray_15_14_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_14_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_14_MPORT_addr = replace_set;
  assign dataArray_15_14_MPORT_mask = _GEN_2032 & _GEN_1581;
  assign dataArray_15_14_MPORT_en = _T_6 & _off_T;
  assign dataArray_15_15_cachedata_MPORT_en = dataArray_15_15_cachedata_MPORT_en_pipe_0;
  assign dataArray_15_15_cachedata_MPORT_addr = dataArray_15_15_cachedata_MPORT_addr_pipe_0;
  assign dataArray_15_15_cachedata_MPORT_data = dataArray_15_15[dataArray_15_15_cachedata_MPORT_addr]; // @[cache.scala 30:33]
  assign dataArray_15_15_MPORT_data = to_sram_r_bits_data;
  assign dataArray_15_15_MPORT_addr = replace_set;
  assign dataArray_15_15_MPORT_mask = _GEN_2032 & _GEN_1583;
  assign dataArray_15_15_MPORT_en = _T_6 & _off_T;
  assign from_IFU_ready = 3'h0 == state_cache; // @[Mux.scala 81:61]
  assign to_IFU_valid = 3'h1 == state_cache; // @[Mux.scala 81:61]
  assign to_IFU_bits_data = hit ? _GEN_1551 : 32'h13; // @[cache.scala 108:28]
  assign to_sram_ar_valid = 3'h2 == state_cache; // @[Mux.scala 81:61]
  assign to_sram_ar_bits_addr = _to_sram_ar_bits_addr_T_3[31:0]; // @[cache.scala 91:27]
  assign to_sram_ar_bits_len = {{4'd0}, _to_sram_ar_bits_len_T_1}; // @[cache.scala 93:27]
  assign to_sram_r_ready = 3'h3 == state_cache; // @[Mux.scala 81:61]
  always @(posedge clock) begin
    if (dataArray_0_0_MPORT_en & dataArray_0_0_MPORT_mask) begin
      dataArray_0_0[dataArray_0_0_MPORT_addr] <= dataArray_0_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_1_MPORT_en & dataArray_0_1_MPORT_mask) begin
      dataArray_0_1[dataArray_0_1_MPORT_addr] <= dataArray_0_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_2_MPORT_en & dataArray_0_2_MPORT_mask) begin
      dataArray_0_2[dataArray_0_2_MPORT_addr] <= dataArray_0_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_3_MPORT_en & dataArray_0_3_MPORT_mask) begin
      dataArray_0_3[dataArray_0_3_MPORT_addr] <= dataArray_0_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_4_MPORT_en & dataArray_0_4_MPORT_mask) begin
      dataArray_0_4[dataArray_0_4_MPORT_addr] <= dataArray_0_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_5_MPORT_en & dataArray_0_5_MPORT_mask) begin
      dataArray_0_5[dataArray_0_5_MPORT_addr] <= dataArray_0_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_6_MPORT_en & dataArray_0_6_MPORT_mask) begin
      dataArray_0_6[dataArray_0_6_MPORT_addr] <= dataArray_0_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_7_MPORT_en & dataArray_0_7_MPORT_mask) begin
      dataArray_0_7[dataArray_0_7_MPORT_addr] <= dataArray_0_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_8_MPORT_en & dataArray_0_8_MPORT_mask) begin
      dataArray_0_8[dataArray_0_8_MPORT_addr] <= dataArray_0_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_9_MPORT_en & dataArray_0_9_MPORT_mask) begin
      dataArray_0_9[dataArray_0_9_MPORT_addr] <= dataArray_0_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_10_MPORT_en & dataArray_0_10_MPORT_mask) begin
      dataArray_0_10[dataArray_0_10_MPORT_addr] <= dataArray_0_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_11_MPORT_en & dataArray_0_11_MPORT_mask) begin
      dataArray_0_11[dataArray_0_11_MPORT_addr] <= dataArray_0_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_12_MPORT_en & dataArray_0_12_MPORT_mask) begin
      dataArray_0_12[dataArray_0_12_MPORT_addr] <= dataArray_0_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_13_MPORT_en & dataArray_0_13_MPORT_mask) begin
      dataArray_0_13[dataArray_0_13_MPORT_addr] <= dataArray_0_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_14_MPORT_en & dataArray_0_14_MPORT_mask) begin
      dataArray_0_14[dataArray_0_14_MPORT_addr] <= dataArray_0_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_0_15_MPORT_en & dataArray_0_15_MPORT_mask) begin
      dataArray_0_15[dataArray_0_15_MPORT_addr] <= dataArray_0_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_0_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_0_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_0_MPORT_en & dataArray_1_0_MPORT_mask) begin
      dataArray_1_0[dataArray_1_0_MPORT_addr] <= dataArray_1_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_1_MPORT_en & dataArray_1_1_MPORT_mask) begin
      dataArray_1_1[dataArray_1_1_MPORT_addr] <= dataArray_1_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_2_MPORT_en & dataArray_1_2_MPORT_mask) begin
      dataArray_1_2[dataArray_1_2_MPORT_addr] <= dataArray_1_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_3_MPORT_en & dataArray_1_3_MPORT_mask) begin
      dataArray_1_3[dataArray_1_3_MPORT_addr] <= dataArray_1_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_4_MPORT_en & dataArray_1_4_MPORT_mask) begin
      dataArray_1_4[dataArray_1_4_MPORT_addr] <= dataArray_1_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_5_MPORT_en & dataArray_1_5_MPORT_mask) begin
      dataArray_1_5[dataArray_1_5_MPORT_addr] <= dataArray_1_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_6_MPORT_en & dataArray_1_6_MPORT_mask) begin
      dataArray_1_6[dataArray_1_6_MPORT_addr] <= dataArray_1_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_7_MPORT_en & dataArray_1_7_MPORT_mask) begin
      dataArray_1_7[dataArray_1_7_MPORT_addr] <= dataArray_1_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_8_MPORT_en & dataArray_1_8_MPORT_mask) begin
      dataArray_1_8[dataArray_1_8_MPORT_addr] <= dataArray_1_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_9_MPORT_en & dataArray_1_9_MPORT_mask) begin
      dataArray_1_9[dataArray_1_9_MPORT_addr] <= dataArray_1_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_10_MPORT_en & dataArray_1_10_MPORT_mask) begin
      dataArray_1_10[dataArray_1_10_MPORT_addr] <= dataArray_1_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_11_MPORT_en & dataArray_1_11_MPORT_mask) begin
      dataArray_1_11[dataArray_1_11_MPORT_addr] <= dataArray_1_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_12_MPORT_en & dataArray_1_12_MPORT_mask) begin
      dataArray_1_12[dataArray_1_12_MPORT_addr] <= dataArray_1_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_13_MPORT_en & dataArray_1_13_MPORT_mask) begin
      dataArray_1_13[dataArray_1_13_MPORT_addr] <= dataArray_1_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_14_MPORT_en & dataArray_1_14_MPORT_mask) begin
      dataArray_1_14[dataArray_1_14_MPORT_addr] <= dataArray_1_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_1_15_MPORT_en & dataArray_1_15_MPORT_mask) begin
      dataArray_1_15[dataArray_1_15_MPORT_addr] <= dataArray_1_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_1_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_1_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_0_MPORT_en & dataArray_2_0_MPORT_mask) begin
      dataArray_2_0[dataArray_2_0_MPORT_addr] <= dataArray_2_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_1_MPORT_en & dataArray_2_1_MPORT_mask) begin
      dataArray_2_1[dataArray_2_1_MPORT_addr] <= dataArray_2_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_2_MPORT_en & dataArray_2_2_MPORT_mask) begin
      dataArray_2_2[dataArray_2_2_MPORT_addr] <= dataArray_2_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_3_MPORT_en & dataArray_2_3_MPORT_mask) begin
      dataArray_2_3[dataArray_2_3_MPORT_addr] <= dataArray_2_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_4_MPORT_en & dataArray_2_4_MPORT_mask) begin
      dataArray_2_4[dataArray_2_4_MPORT_addr] <= dataArray_2_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_5_MPORT_en & dataArray_2_5_MPORT_mask) begin
      dataArray_2_5[dataArray_2_5_MPORT_addr] <= dataArray_2_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_6_MPORT_en & dataArray_2_6_MPORT_mask) begin
      dataArray_2_6[dataArray_2_6_MPORT_addr] <= dataArray_2_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_7_MPORT_en & dataArray_2_7_MPORT_mask) begin
      dataArray_2_7[dataArray_2_7_MPORT_addr] <= dataArray_2_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_8_MPORT_en & dataArray_2_8_MPORT_mask) begin
      dataArray_2_8[dataArray_2_8_MPORT_addr] <= dataArray_2_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_9_MPORT_en & dataArray_2_9_MPORT_mask) begin
      dataArray_2_9[dataArray_2_9_MPORT_addr] <= dataArray_2_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_10_MPORT_en & dataArray_2_10_MPORT_mask) begin
      dataArray_2_10[dataArray_2_10_MPORT_addr] <= dataArray_2_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_11_MPORT_en & dataArray_2_11_MPORT_mask) begin
      dataArray_2_11[dataArray_2_11_MPORT_addr] <= dataArray_2_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_12_MPORT_en & dataArray_2_12_MPORT_mask) begin
      dataArray_2_12[dataArray_2_12_MPORT_addr] <= dataArray_2_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_13_MPORT_en & dataArray_2_13_MPORT_mask) begin
      dataArray_2_13[dataArray_2_13_MPORT_addr] <= dataArray_2_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_14_MPORT_en & dataArray_2_14_MPORT_mask) begin
      dataArray_2_14[dataArray_2_14_MPORT_addr] <= dataArray_2_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_2_15_MPORT_en & dataArray_2_15_MPORT_mask) begin
      dataArray_2_15[dataArray_2_15_MPORT_addr] <= dataArray_2_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_2_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_2_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_0_MPORT_en & dataArray_3_0_MPORT_mask) begin
      dataArray_3_0[dataArray_3_0_MPORT_addr] <= dataArray_3_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_1_MPORT_en & dataArray_3_1_MPORT_mask) begin
      dataArray_3_1[dataArray_3_1_MPORT_addr] <= dataArray_3_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_2_MPORT_en & dataArray_3_2_MPORT_mask) begin
      dataArray_3_2[dataArray_3_2_MPORT_addr] <= dataArray_3_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_3_MPORT_en & dataArray_3_3_MPORT_mask) begin
      dataArray_3_3[dataArray_3_3_MPORT_addr] <= dataArray_3_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_4_MPORT_en & dataArray_3_4_MPORT_mask) begin
      dataArray_3_4[dataArray_3_4_MPORT_addr] <= dataArray_3_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_5_MPORT_en & dataArray_3_5_MPORT_mask) begin
      dataArray_3_5[dataArray_3_5_MPORT_addr] <= dataArray_3_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_6_MPORT_en & dataArray_3_6_MPORT_mask) begin
      dataArray_3_6[dataArray_3_6_MPORT_addr] <= dataArray_3_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_7_MPORT_en & dataArray_3_7_MPORT_mask) begin
      dataArray_3_7[dataArray_3_7_MPORT_addr] <= dataArray_3_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_8_MPORT_en & dataArray_3_8_MPORT_mask) begin
      dataArray_3_8[dataArray_3_8_MPORT_addr] <= dataArray_3_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_9_MPORT_en & dataArray_3_9_MPORT_mask) begin
      dataArray_3_9[dataArray_3_9_MPORT_addr] <= dataArray_3_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_10_MPORT_en & dataArray_3_10_MPORT_mask) begin
      dataArray_3_10[dataArray_3_10_MPORT_addr] <= dataArray_3_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_11_MPORT_en & dataArray_3_11_MPORT_mask) begin
      dataArray_3_11[dataArray_3_11_MPORT_addr] <= dataArray_3_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_12_MPORT_en & dataArray_3_12_MPORT_mask) begin
      dataArray_3_12[dataArray_3_12_MPORT_addr] <= dataArray_3_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_13_MPORT_en & dataArray_3_13_MPORT_mask) begin
      dataArray_3_13[dataArray_3_13_MPORT_addr] <= dataArray_3_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_14_MPORT_en & dataArray_3_14_MPORT_mask) begin
      dataArray_3_14[dataArray_3_14_MPORT_addr] <= dataArray_3_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_3_15_MPORT_en & dataArray_3_15_MPORT_mask) begin
      dataArray_3_15[dataArray_3_15_MPORT_addr] <= dataArray_3_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_3_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_3_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_0_MPORT_en & dataArray_4_0_MPORT_mask) begin
      dataArray_4_0[dataArray_4_0_MPORT_addr] <= dataArray_4_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_1_MPORT_en & dataArray_4_1_MPORT_mask) begin
      dataArray_4_1[dataArray_4_1_MPORT_addr] <= dataArray_4_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_2_MPORT_en & dataArray_4_2_MPORT_mask) begin
      dataArray_4_2[dataArray_4_2_MPORT_addr] <= dataArray_4_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_3_MPORT_en & dataArray_4_3_MPORT_mask) begin
      dataArray_4_3[dataArray_4_3_MPORT_addr] <= dataArray_4_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_4_MPORT_en & dataArray_4_4_MPORT_mask) begin
      dataArray_4_4[dataArray_4_4_MPORT_addr] <= dataArray_4_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_5_MPORT_en & dataArray_4_5_MPORT_mask) begin
      dataArray_4_5[dataArray_4_5_MPORT_addr] <= dataArray_4_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_6_MPORT_en & dataArray_4_6_MPORT_mask) begin
      dataArray_4_6[dataArray_4_6_MPORT_addr] <= dataArray_4_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_7_MPORT_en & dataArray_4_7_MPORT_mask) begin
      dataArray_4_7[dataArray_4_7_MPORT_addr] <= dataArray_4_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_8_MPORT_en & dataArray_4_8_MPORT_mask) begin
      dataArray_4_8[dataArray_4_8_MPORT_addr] <= dataArray_4_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_9_MPORT_en & dataArray_4_9_MPORT_mask) begin
      dataArray_4_9[dataArray_4_9_MPORT_addr] <= dataArray_4_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_10_MPORT_en & dataArray_4_10_MPORT_mask) begin
      dataArray_4_10[dataArray_4_10_MPORT_addr] <= dataArray_4_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_11_MPORT_en & dataArray_4_11_MPORT_mask) begin
      dataArray_4_11[dataArray_4_11_MPORT_addr] <= dataArray_4_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_12_MPORT_en & dataArray_4_12_MPORT_mask) begin
      dataArray_4_12[dataArray_4_12_MPORT_addr] <= dataArray_4_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_13_MPORT_en & dataArray_4_13_MPORT_mask) begin
      dataArray_4_13[dataArray_4_13_MPORT_addr] <= dataArray_4_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_14_MPORT_en & dataArray_4_14_MPORT_mask) begin
      dataArray_4_14[dataArray_4_14_MPORT_addr] <= dataArray_4_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_4_15_MPORT_en & dataArray_4_15_MPORT_mask) begin
      dataArray_4_15[dataArray_4_15_MPORT_addr] <= dataArray_4_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_4_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_4_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_0_MPORT_en & dataArray_5_0_MPORT_mask) begin
      dataArray_5_0[dataArray_5_0_MPORT_addr] <= dataArray_5_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_1_MPORT_en & dataArray_5_1_MPORT_mask) begin
      dataArray_5_1[dataArray_5_1_MPORT_addr] <= dataArray_5_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_2_MPORT_en & dataArray_5_2_MPORT_mask) begin
      dataArray_5_2[dataArray_5_2_MPORT_addr] <= dataArray_5_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_3_MPORT_en & dataArray_5_3_MPORT_mask) begin
      dataArray_5_3[dataArray_5_3_MPORT_addr] <= dataArray_5_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_4_MPORT_en & dataArray_5_4_MPORT_mask) begin
      dataArray_5_4[dataArray_5_4_MPORT_addr] <= dataArray_5_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_5_MPORT_en & dataArray_5_5_MPORT_mask) begin
      dataArray_5_5[dataArray_5_5_MPORT_addr] <= dataArray_5_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_6_MPORT_en & dataArray_5_6_MPORT_mask) begin
      dataArray_5_6[dataArray_5_6_MPORT_addr] <= dataArray_5_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_7_MPORT_en & dataArray_5_7_MPORT_mask) begin
      dataArray_5_7[dataArray_5_7_MPORT_addr] <= dataArray_5_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_8_MPORT_en & dataArray_5_8_MPORT_mask) begin
      dataArray_5_8[dataArray_5_8_MPORT_addr] <= dataArray_5_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_9_MPORT_en & dataArray_5_9_MPORT_mask) begin
      dataArray_5_9[dataArray_5_9_MPORT_addr] <= dataArray_5_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_10_MPORT_en & dataArray_5_10_MPORT_mask) begin
      dataArray_5_10[dataArray_5_10_MPORT_addr] <= dataArray_5_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_11_MPORT_en & dataArray_5_11_MPORT_mask) begin
      dataArray_5_11[dataArray_5_11_MPORT_addr] <= dataArray_5_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_12_MPORT_en & dataArray_5_12_MPORT_mask) begin
      dataArray_5_12[dataArray_5_12_MPORT_addr] <= dataArray_5_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_13_MPORT_en & dataArray_5_13_MPORT_mask) begin
      dataArray_5_13[dataArray_5_13_MPORT_addr] <= dataArray_5_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_14_MPORT_en & dataArray_5_14_MPORT_mask) begin
      dataArray_5_14[dataArray_5_14_MPORT_addr] <= dataArray_5_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_5_15_MPORT_en & dataArray_5_15_MPORT_mask) begin
      dataArray_5_15[dataArray_5_15_MPORT_addr] <= dataArray_5_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_5_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_5_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_0_MPORT_en & dataArray_6_0_MPORT_mask) begin
      dataArray_6_0[dataArray_6_0_MPORT_addr] <= dataArray_6_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_1_MPORT_en & dataArray_6_1_MPORT_mask) begin
      dataArray_6_1[dataArray_6_1_MPORT_addr] <= dataArray_6_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_2_MPORT_en & dataArray_6_2_MPORT_mask) begin
      dataArray_6_2[dataArray_6_2_MPORT_addr] <= dataArray_6_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_3_MPORT_en & dataArray_6_3_MPORT_mask) begin
      dataArray_6_3[dataArray_6_3_MPORT_addr] <= dataArray_6_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_4_MPORT_en & dataArray_6_4_MPORT_mask) begin
      dataArray_6_4[dataArray_6_4_MPORT_addr] <= dataArray_6_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_5_MPORT_en & dataArray_6_5_MPORT_mask) begin
      dataArray_6_5[dataArray_6_5_MPORT_addr] <= dataArray_6_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_6_MPORT_en & dataArray_6_6_MPORT_mask) begin
      dataArray_6_6[dataArray_6_6_MPORT_addr] <= dataArray_6_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_7_MPORT_en & dataArray_6_7_MPORT_mask) begin
      dataArray_6_7[dataArray_6_7_MPORT_addr] <= dataArray_6_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_8_MPORT_en & dataArray_6_8_MPORT_mask) begin
      dataArray_6_8[dataArray_6_8_MPORT_addr] <= dataArray_6_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_9_MPORT_en & dataArray_6_9_MPORT_mask) begin
      dataArray_6_9[dataArray_6_9_MPORT_addr] <= dataArray_6_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_10_MPORT_en & dataArray_6_10_MPORT_mask) begin
      dataArray_6_10[dataArray_6_10_MPORT_addr] <= dataArray_6_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_11_MPORT_en & dataArray_6_11_MPORT_mask) begin
      dataArray_6_11[dataArray_6_11_MPORT_addr] <= dataArray_6_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_12_MPORT_en & dataArray_6_12_MPORT_mask) begin
      dataArray_6_12[dataArray_6_12_MPORT_addr] <= dataArray_6_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_13_MPORT_en & dataArray_6_13_MPORT_mask) begin
      dataArray_6_13[dataArray_6_13_MPORT_addr] <= dataArray_6_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_14_MPORT_en & dataArray_6_14_MPORT_mask) begin
      dataArray_6_14[dataArray_6_14_MPORT_addr] <= dataArray_6_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_6_15_MPORT_en & dataArray_6_15_MPORT_mask) begin
      dataArray_6_15[dataArray_6_15_MPORT_addr] <= dataArray_6_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_6_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_6_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_0_MPORT_en & dataArray_7_0_MPORT_mask) begin
      dataArray_7_0[dataArray_7_0_MPORT_addr] <= dataArray_7_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_1_MPORT_en & dataArray_7_1_MPORT_mask) begin
      dataArray_7_1[dataArray_7_1_MPORT_addr] <= dataArray_7_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_2_MPORT_en & dataArray_7_2_MPORT_mask) begin
      dataArray_7_2[dataArray_7_2_MPORT_addr] <= dataArray_7_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_3_MPORT_en & dataArray_7_3_MPORT_mask) begin
      dataArray_7_3[dataArray_7_3_MPORT_addr] <= dataArray_7_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_4_MPORT_en & dataArray_7_4_MPORT_mask) begin
      dataArray_7_4[dataArray_7_4_MPORT_addr] <= dataArray_7_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_5_MPORT_en & dataArray_7_5_MPORT_mask) begin
      dataArray_7_5[dataArray_7_5_MPORT_addr] <= dataArray_7_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_6_MPORT_en & dataArray_7_6_MPORT_mask) begin
      dataArray_7_6[dataArray_7_6_MPORT_addr] <= dataArray_7_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_7_MPORT_en & dataArray_7_7_MPORT_mask) begin
      dataArray_7_7[dataArray_7_7_MPORT_addr] <= dataArray_7_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_8_MPORT_en & dataArray_7_8_MPORT_mask) begin
      dataArray_7_8[dataArray_7_8_MPORT_addr] <= dataArray_7_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_9_MPORT_en & dataArray_7_9_MPORT_mask) begin
      dataArray_7_9[dataArray_7_9_MPORT_addr] <= dataArray_7_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_10_MPORT_en & dataArray_7_10_MPORT_mask) begin
      dataArray_7_10[dataArray_7_10_MPORT_addr] <= dataArray_7_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_11_MPORT_en & dataArray_7_11_MPORT_mask) begin
      dataArray_7_11[dataArray_7_11_MPORT_addr] <= dataArray_7_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_12_MPORT_en & dataArray_7_12_MPORT_mask) begin
      dataArray_7_12[dataArray_7_12_MPORT_addr] <= dataArray_7_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_13_MPORT_en & dataArray_7_13_MPORT_mask) begin
      dataArray_7_13[dataArray_7_13_MPORT_addr] <= dataArray_7_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_14_MPORT_en & dataArray_7_14_MPORT_mask) begin
      dataArray_7_14[dataArray_7_14_MPORT_addr] <= dataArray_7_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_7_15_MPORT_en & dataArray_7_15_MPORT_mask) begin
      dataArray_7_15[dataArray_7_15_MPORT_addr] <= dataArray_7_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_7_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_7_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_0_MPORT_en & dataArray_8_0_MPORT_mask) begin
      dataArray_8_0[dataArray_8_0_MPORT_addr] <= dataArray_8_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_1_MPORT_en & dataArray_8_1_MPORT_mask) begin
      dataArray_8_1[dataArray_8_1_MPORT_addr] <= dataArray_8_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_2_MPORT_en & dataArray_8_2_MPORT_mask) begin
      dataArray_8_2[dataArray_8_2_MPORT_addr] <= dataArray_8_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_3_MPORT_en & dataArray_8_3_MPORT_mask) begin
      dataArray_8_3[dataArray_8_3_MPORT_addr] <= dataArray_8_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_4_MPORT_en & dataArray_8_4_MPORT_mask) begin
      dataArray_8_4[dataArray_8_4_MPORT_addr] <= dataArray_8_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_5_MPORT_en & dataArray_8_5_MPORT_mask) begin
      dataArray_8_5[dataArray_8_5_MPORT_addr] <= dataArray_8_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_6_MPORT_en & dataArray_8_6_MPORT_mask) begin
      dataArray_8_6[dataArray_8_6_MPORT_addr] <= dataArray_8_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_7_MPORT_en & dataArray_8_7_MPORT_mask) begin
      dataArray_8_7[dataArray_8_7_MPORT_addr] <= dataArray_8_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_8_MPORT_en & dataArray_8_8_MPORT_mask) begin
      dataArray_8_8[dataArray_8_8_MPORT_addr] <= dataArray_8_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_9_MPORT_en & dataArray_8_9_MPORT_mask) begin
      dataArray_8_9[dataArray_8_9_MPORT_addr] <= dataArray_8_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_10_MPORT_en & dataArray_8_10_MPORT_mask) begin
      dataArray_8_10[dataArray_8_10_MPORT_addr] <= dataArray_8_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_11_MPORT_en & dataArray_8_11_MPORT_mask) begin
      dataArray_8_11[dataArray_8_11_MPORT_addr] <= dataArray_8_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_12_MPORT_en & dataArray_8_12_MPORT_mask) begin
      dataArray_8_12[dataArray_8_12_MPORT_addr] <= dataArray_8_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_13_MPORT_en & dataArray_8_13_MPORT_mask) begin
      dataArray_8_13[dataArray_8_13_MPORT_addr] <= dataArray_8_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_14_MPORT_en & dataArray_8_14_MPORT_mask) begin
      dataArray_8_14[dataArray_8_14_MPORT_addr] <= dataArray_8_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_8_15_MPORT_en & dataArray_8_15_MPORT_mask) begin
      dataArray_8_15[dataArray_8_15_MPORT_addr] <= dataArray_8_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_8_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_8_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_0_MPORT_en & dataArray_9_0_MPORT_mask) begin
      dataArray_9_0[dataArray_9_0_MPORT_addr] <= dataArray_9_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_1_MPORT_en & dataArray_9_1_MPORT_mask) begin
      dataArray_9_1[dataArray_9_1_MPORT_addr] <= dataArray_9_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_2_MPORT_en & dataArray_9_2_MPORT_mask) begin
      dataArray_9_2[dataArray_9_2_MPORT_addr] <= dataArray_9_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_3_MPORT_en & dataArray_9_3_MPORT_mask) begin
      dataArray_9_3[dataArray_9_3_MPORT_addr] <= dataArray_9_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_4_MPORT_en & dataArray_9_4_MPORT_mask) begin
      dataArray_9_4[dataArray_9_4_MPORT_addr] <= dataArray_9_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_5_MPORT_en & dataArray_9_5_MPORT_mask) begin
      dataArray_9_5[dataArray_9_5_MPORT_addr] <= dataArray_9_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_6_MPORT_en & dataArray_9_6_MPORT_mask) begin
      dataArray_9_6[dataArray_9_6_MPORT_addr] <= dataArray_9_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_7_MPORT_en & dataArray_9_7_MPORT_mask) begin
      dataArray_9_7[dataArray_9_7_MPORT_addr] <= dataArray_9_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_8_MPORT_en & dataArray_9_8_MPORT_mask) begin
      dataArray_9_8[dataArray_9_8_MPORT_addr] <= dataArray_9_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_9_MPORT_en & dataArray_9_9_MPORT_mask) begin
      dataArray_9_9[dataArray_9_9_MPORT_addr] <= dataArray_9_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_10_MPORT_en & dataArray_9_10_MPORT_mask) begin
      dataArray_9_10[dataArray_9_10_MPORT_addr] <= dataArray_9_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_11_MPORT_en & dataArray_9_11_MPORT_mask) begin
      dataArray_9_11[dataArray_9_11_MPORT_addr] <= dataArray_9_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_12_MPORT_en & dataArray_9_12_MPORT_mask) begin
      dataArray_9_12[dataArray_9_12_MPORT_addr] <= dataArray_9_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_13_MPORT_en & dataArray_9_13_MPORT_mask) begin
      dataArray_9_13[dataArray_9_13_MPORT_addr] <= dataArray_9_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_14_MPORT_en & dataArray_9_14_MPORT_mask) begin
      dataArray_9_14[dataArray_9_14_MPORT_addr] <= dataArray_9_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_9_15_MPORT_en & dataArray_9_15_MPORT_mask) begin
      dataArray_9_15[dataArray_9_15_MPORT_addr] <= dataArray_9_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_9_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_9_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_0_MPORT_en & dataArray_10_0_MPORT_mask) begin
      dataArray_10_0[dataArray_10_0_MPORT_addr] <= dataArray_10_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_1_MPORT_en & dataArray_10_1_MPORT_mask) begin
      dataArray_10_1[dataArray_10_1_MPORT_addr] <= dataArray_10_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_2_MPORT_en & dataArray_10_2_MPORT_mask) begin
      dataArray_10_2[dataArray_10_2_MPORT_addr] <= dataArray_10_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_3_MPORT_en & dataArray_10_3_MPORT_mask) begin
      dataArray_10_3[dataArray_10_3_MPORT_addr] <= dataArray_10_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_4_MPORT_en & dataArray_10_4_MPORT_mask) begin
      dataArray_10_4[dataArray_10_4_MPORT_addr] <= dataArray_10_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_5_MPORT_en & dataArray_10_5_MPORT_mask) begin
      dataArray_10_5[dataArray_10_5_MPORT_addr] <= dataArray_10_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_6_MPORT_en & dataArray_10_6_MPORT_mask) begin
      dataArray_10_6[dataArray_10_6_MPORT_addr] <= dataArray_10_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_7_MPORT_en & dataArray_10_7_MPORT_mask) begin
      dataArray_10_7[dataArray_10_7_MPORT_addr] <= dataArray_10_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_8_MPORT_en & dataArray_10_8_MPORT_mask) begin
      dataArray_10_8[dataArray_10_8_MPORT_addr] <= dataArray_10_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_9_MPORT_en & dataArray_10_9_MPORT_mask) begin
      dataArray_10_9[dataArray_10_9_MPORT_addr] <= dataArray_10_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_10_MPORT_en & dataArray_10_10_MPORT_mask) begin
      dataArray_10_10[dataArray_10_10_MPORT_addr] <= dataArray_10_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_11_MPORT_en & dataArray_10_11_MPORT_mask) begin
      dataArray_10_11[dataArray_10_11_MPORT_addr] <= dataArray_10_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_12_MPORT_en & dataArray_10_12_MPORT_mask) begin
      dataArray_10_12[dataArray_10_12_MPORT_addr] <= dataArray_10_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_13_MPORT_en & dataArray_10_13_MPORT_mask) begin
      dataArray_10_13[dataArray_10_13_MPORT_addr] <= dataArray_10_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_14_MPORT_en & dataArray_10_14_MPORT_mask) begin
      dataArray_10_14[dataArray_10_14_MPORT_addr] <= dataArray_10_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_10_15_MPORT_en & dataArray_10_15_MPORT_mask) begin
      dataArray_10_15[dataArray_10_15_MPORT_addr] <= dataArray_10_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_10_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_10_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_0_MPORT_en & dataArray_11_0_MPORT_mask) begin
      dataArray_11_0[dataArray_11_0_MPORT_addr] <= dataArray_11_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_1_MPORT_en & dataArray_11_1_MPORT_mask) begin
      dataArray_11_1[dataArray_11_1_MPORT_addr] <= dataArray_11_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_2_MPORT_en & dataArray_11_2_MPORT_mask) begin
      dataArray_11_2[dataArray_11_2_MPORT_addr] <= dataArray_11_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_3_MPORT_en & dataArray_11_3_MPORT_mask) begin
      dataArray_11_3[dataArray_11_3_MPORT_addr] <= dataArray_11_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_4_MPORT_en & dataArray_11_4_MPORT_mask) begin
      dataArray_11_4[dataArray_11_4_MPORT_addr] <= dataArray_11_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_5_MPORT_en & dataArray_11_5_MPORT_mask) begin
      dataArray_11_5[dataArray_11_5_MPORT_addr] <= dataArray_11_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_6_MPORT_en & dataArray_11_6_MPORT_mask) begin
      dataArray_11_6[dataArray_11_6_MPORT_addr] <= dataArray_11_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_7_MPORT_en & dataArray_11_7_MPORT_mask) begin
      dataArray_11_7[dataArray_11_7_MPORT_addr] <= dataArray_11_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_8_MPORT_en & dataArray_11_8_MPORT_mask) begin
      dataArray_11_8[dataArray_11_8_MPORT_addr] <= dataArray_11_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_9_MPORT_en & dataArray_11_9_MPORT_mask) begin
      dataArray_11_9[dataArray_11_9_MPORT_addr] <= dataArray_11_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_10_MPORT_en & dataArray_11_10_MPORT_mask) begin
      dataArray_11_10[dataArray_11_10_MPORT_addr] <= dataArray_11_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_11_MPORT_en & dataArray_11_11_MPORT_mask) begin
      dataArray_11_11[dataArray_11_11_MPORT_addr] <= dataArray_11_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_12_MPORT_en & dataArray_11_12_MPORT_mask) begin
      dataArray_11_12[dataArray_11_12_MPORT_addr] <= dataArray_11_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_13_MPORT_en & dataArray_11_13_MPORT_mask) begin
      dataArray_11_13[dataArray_11_13_MPORT_addr] <= dataArray_11_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_14_MPORT_en & dataArray_11_14_MPORT_mask) begin
      dataArray_11_14[dataArray_11_14_MPORT_addr] <= dataArray_11_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_11_15_MPORT_en & dataArray_11_15_MPORT_mask) begin
      dataArray_11_15[dataArray_11_15_MPORT_addr] <= dataArray_11_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_11_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_11_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_0_MPORT_en & dataArray_12_0_MPORT_mask) begin
      dataArray_12_0[dataArray_12_0_MPORT_addr] <= dataArray_12_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_1_MPORT_en & dataArray_12_1_MPORT_mask) begin
      dataArray_12_1[dataArray_12_1_MPORT_addr] <= dataArray_12_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_2_MPORT_en & dataArray_12_2_MPORT_mask) begin
      dataArray_12_2[dataArray_12_2_MPORT_addr] <= dataArray_12_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_3_MPORT_en & dataArray_12_3_MPORT_mask) begin
      dataArray_12_3[dataArray_12_3_MPORT_addr] <= dataArray_12_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_4_MPORT_en & dataArray_12_4_MPORT_mask) begin
      dataArray_12_4[dataArray_12_4_MPORT_addr] <= dataArray_12_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_5_MPORT_en & dataArray_12_5_MPORT_mask) begin
      dataArray_12_5[dataArray_12_5_MPORT_addr] <= dataArray_12_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_6_MPORT_en & dataArray_12_6_MPORT_mask) begin
      dataArray_12_6[dataArray_12_6_MPORT_addr] <= dataArray_12_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_7_MPORT_en & dataArray_12_7_MPORT_mask) begin
      dataArray_12_7[dataArray_12_7_MPORT_addr] <= dataArray_12_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_8_MPORT_en & dataArray_12_8_MPORT_mask) begin
      dataArray_12_8[dataArray_12_8_MPORT_addr] <= dataArray_12_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_9_MPORT_en & dataArray_12_9_MPORT_mask) begin
      dataArray_12_9[dataArray_12_9_MPORT_addr] <= dataArray_12_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_10_MPORT_en & dataArray_12_10_MPORT_mask) begin
      dataArray_12_10[dataArray_12_10_MPORT_addr] <= dataArray_12_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_11_MPORT_en & dataArray_12_11_MPORT_mask) begin
      dataArray_12_11[dataArray_12_11_MPORT_addr] <= dataArray_12_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_12_MPORT_en & dataArray_12_12_MPORT_mask) begin
      dataArray_12_12[dataArray_12_12_MPORT_addr] <= dataArray_12_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_13_MPORT_en & dataArray_12_13_MPORT_mask) begin
      dataArray_12_13[dataArray_12_13_MPORT_addr] <= dataArray_12_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_14_MPORT_en & dataArray_12_14_MPORT_mask) begin
      dataArray_12_14[dataArray_12_14_MPORT_addr] <= dataArray_12_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_12_15_MPORT_en & dataArray_12_15_MPORT_mask) begin
      dataArray_12_15[dataArray_12_15_MPORT_addr] <= dataArray_12_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_12_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_12_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_0_MPORT_en & dataArray_13_0_MPORT_mask) begin
      dataArray_13_0[dataArray_13_0_MPORT_addr] <= dataArray_13_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_1_MPORT_en & dataArray_13_1_MPORT_mask) begin
      dataArray_13_1[dataArray_13_1_MPORT_addr] <= dataArray_13_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_2_MPORT_en & dataArray_13_2_MPORT_mask) begin
      dataArray_13_2[dataArray_13_2_MPORT_addr] <= dataArray_13_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_3_MPORT_en & dataArray_13_3_MPORT_mask) begin
      dataArray_13_3[dataArray_13_3_MPORT_addr] <= dataArray_13_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_4_MPORT_en & dataArray_13_4_MPORT_mask) begin
      dataArray_13_4[dataArray_13_4_MPORT_addr] <= dataArray_13_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_5_MPORT_en & dataArray_13_5_MPORT_mask) begin
      dataArray_13_5[dataArray_13_5_MPORT_addr] <= dataArray_13_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_6_MPORT_en & dataArray_13_6_MPORT_mask) begin
      dataArray_13_6[dataArray_13_6_MPORT_addr] <= dataArray_13_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_7_MPORT_en & dataArray_13_7_MPORT_mask) begin
      dataArray_13_7[dataArray_13_7_MPORT_addr] <= dataArray_13_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_8_MPORT_en & dataArray_13_8_MPORT_mask) begin
      dataArray_13_8[dataArray_13_8_MPORT_addr] <= dataArray_13_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_9_MPORT_en & dataArray_13_9_MPORT_mask) begin
      dataArray_13_9[dataArray_13_9_MPORT_addr] <= dataArray_13_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_10_MPORT_en & dataArray_13_10_MPORT_mask) begin
      dataArray_13_10[dataArray_13_10_MPORT_addr] <= dataArray_13_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_11_MPORT_en & dataArray_13_11_MPORT_mask) begin
      dataArray_13_11[dataArray_13_11_MPORT_addr] <= dataArray_13_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_12_MPORT_en & dataArray_13_12_MPORT_mask) begin
      dataArray_13_12[dataArray_13_12_MPORT_addr] <= dataArray_13_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_13_MPORT_en & dataArray_13_13_MPORT_mask) begin
      dataArray_13_13[dataArray_13_13_MPORT_addr] <= dataArray_13_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_14_MPORT_en & dataArray_13_14_MPORT_mask) begin
      dataArray_13_14[dataArray_13_14_MPORT_addr] <= dataArray_13_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_13_15_MPORT_en & dataArray_13_15_MPORT_mask) begin
      dataArray_13_15[dataArray_13_15_MPORT_addr] <= dataArray_13_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_13_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_13_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_0_MPORT_en & dataArray_14_0_MPORT_mask) begin
      dataArray_14_0[dataArray_14_0_MPORT_addr] <= dataArray_14_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_1_MPORT_en & dataArray_14_1_MPORT_mask) begin
      dataArray_14_1[dataArray_14_1_MPORT_addr] <= dataArray_14_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_2_MPORT_en & dataArray_14_2_MPORT_mask) begin
      dataArray_14_2[dataArray_14_2_MPORT_addr] <= dataArray_14_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_3_MPORT_en & dataArray_14_3_MPORT_mask) begin
      dataArray_14_3[dataArray_14_3_MPORT_addr] <= dataArray_14_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_4_MPORT_en & dataArray_14_4_MPORT_mask) begin
      dataArray_14_4[dataArray_14_4_MPORT_addr] <= dataArray_14_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_5_MPORT_en & dataArray_14_5_MPORT_mask) begin
      dataArray_14_5[dataArray_14_5_MPORT_addr] <= dataArray_14_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_6_MPORT_en & dataArray_14_6_MPORT_mask) begin
      dataArray_14_6[dataArray_14_6_MPORT_addr] <= dataArray_14_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_7_MPORT_en & dataArray_14_7_MPORT_mask) begin
      dataArray_14_7[dataArray_14_7_MPORT_addr] <= dataArray_14_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_8_MPORT_en & dataArray_14_8_MPORT_mask) begin
      dataArray_14_8[dataArray_14_8_MPORT_addr] <= dataArray_14_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_9_MPORT_en & dataArray_14_9_MPORT_mask) begin
      dataArray_14_9[dataArray_14_9_MPORT_addr] <= dataArray_14_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_10_MPORT_en & dataArray_14_10_MPORT_mask) begin
      dataArray_14_10[dataArray_14_10_MPORT_addr] <= dataArray_14_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_11_MPORT_en & dataArray_14_11_MPORT_mask) begin
      dataArray_14_11[dataArray_14_11_MPORT_addr] <= dataArray_14_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_12_MPORT_en & dataArray_14_12_MPORT_mask) begin
      dataArray_14_12[dataArray_14_12_MPORT_addr] <= dataArray_14_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_13_MPORT_en & dataArray_14_13_MPORT_mask) begin
      dataArray_14_13[dataArray_14_13_MPORT_addr] <= dataArray_14_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_14_MPORT_en & dataArray_14_14_MPORT_mask) begin
      dataArray_14_14[dataArray_14_14_MPORT_addr] <= dataArray_14_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_14_15_MPORT_en & dataArray_14_15_MPORT_mask) begin
      dataArray_14_15[dataArray_14_15_MPORT_addr] <= dataArray_14_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_14_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_14_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_0_MPORT_en & dataArray_15_0_MPORT_mask) begin
      dataArray_15_0[dataArray_15_0_MPORT_addr] <= dataArray_15_0_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_0_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_0_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_1_MPORT_en & dataArray_15_1_MPORT_mask) begin
      dataArray_15_1[dataArray_15_1_MPORT_addr] <= dataArray_15_1_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_1_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_1_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_2_MPORT_en & dataArray_15_2_MPORT_mask) begin
      dataArray_15_2[dataArray_15_2_MPORT_addr] <= dataArray_15_2_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_2_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_2_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_3_MPORT_en & dataArray_15_3_MPORT_mask) begin
      dataArray_15_3[dataArray_15_3_MPORT_addr] <= dataArray_15_3_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_3_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_3_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_4_MPORT_en & dataArray_15_4_MPORT_mask) begin
      dataArray_15_4[dataArray_15_4_MPORT_addr] <= dataArray_15_4_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_4_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_4_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_5_MPORT_en & dataArray_15_5_MPORT_mask) begin
      dataArray_15_5[dataArray_15_5_MPORT_addr] <= dataArray_15_5_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_5_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_5_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_6_MPORT_en & dataArray_15_6_MPORT_mask) begin
      dataArray_15_6[dataArray_15_6_MPORT_addr] <= dataArray_15_6_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_6_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_6_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_7_MPORT_en & dataArray_15_7_MPORT_mask) begin
      dataArray_15_7[dataArray_15_7_MPORT_addr] <= dataArray_15_7_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_7_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_7_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_8_MPORT_en & dataArray_15_8_MPORT_mask) begin
      dataArray_15_8[dataArray_15_8_MPORT_addr] <= dataArray_15_8_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_8_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_8_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_9_MPORT_en & dataArray_15_9_MPORT_mask) begin
      dataArray_15_9[dataArray_15_9_MPORT_addr] <= dataArray_15_9_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_9_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_9_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_10_MPORT_en & dataArray_15_10_MPORT_mask) begin
      dataArray_15_10[dataArray_15_10_MPORT_addr] <= dataArray_15_10_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_10_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_10_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_11_MPORT_en & dataArray_15_11_MPORT_mask) begin
      dataArray_15_11[dataArray_15_11_MPORT_addr] <= dataArray_15_11_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_11_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_11_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_12_MPORT_en & dataArray_15_12_MPORT_mask) begin
      dataArray_15_12[dataArray_15_12_MPORT_addr] <= dataArray_15_12_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_12_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_12_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_13_MPORT_en & dataArray_15_13_MPORT_mask) begin
      dataArray_15_13[dataArray_15_13_MPORT_addr] <= dataArray_15_13_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_13_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_13_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_14_MPORT_en & dataArray_15_14_MPORT_mask) begin
      dataArray_15_14[dataArray_15_14_MPORT_addr] <= dataArray_15_14_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_14_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_14_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (dataArray_15_15_MPORT_en & dataArray_15_15_MPORT_mask) begin
      dataArray_15_15[dataArray_15_15_MPORT_addr] <= dataArray_15_15_MPORT_data; // @[cache.scala 30:33]
    end
    dataArray_15_15_cachedata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dataArray_15_15_cachedata_MPORT_addr_pipe_0 <= _GEN_47 == tag;
    end
    if (reset) begin // @[cache.scala 21:30]
      replace_set <= 1'h0; // @[cache.scala 21:30]
    end else if (!(3'h0 == state_cache)) begin // @[cache.scala 49:26]
      if (!(3'h1 == state_cache)) begin // @[cache.scala 49:26]
        if (3'h2 == state_cache) begin // @[cache.scala 49:26]
          replace_set <= random_num; // @[cache.scala 64:25]
        end
      end
    end
    if (reset) begin // @[cache.scala 27:29]
      random_num <= 1'h0; // @[cache.scala 27:29]
    end else begin
      random_num <= random_num + 1'h1; // @[cache.scala 28:16]
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_0 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1552) begin // @[cache.scala 84:50]
          tagArray_0_0 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_1 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1584) begin // @[cache.scala 84:50]
          tagArray_0_1 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_2 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1616) begin // @[cache.scala 84:50]
          tagArray_0_2 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_3 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1648) begin // @[cache.scala 84:50]
          tagArray_0_3 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_4 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1680) begin // @[cache.scala 84:50]
          tagArray_0_4 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_5 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1712) begin // @[cache.scala 84:50]
          tagArray_0_5 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_6 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1744) begin // @[cache.scala 84:50]
          tagArray_0_6 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_7 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1776) begin // @[cache.scala 84:50]
          tagArray_0_7 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_8 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1808) begin // @[cache.scala 84:50]
          tagArray_0_8 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_9 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1840) begin // @[cache.scala 84:50]
          tagArray_0_9 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_10 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1872) begin // @[cache.scala 84:50]
          tagArray_0_10 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_11 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1904) begin // @[cache.scala 84:50]
          tagArray_0_11 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_12 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1936) begin // @[cache.scala 84:50]
          tagArray_0_12 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_13 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_1968) begin // @[cache.scala 84:50]
          tagArray_0_13 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_14 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_2000) begin // @[cache.scala 84:50]
          tagArray_0_14 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_0_15 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (_GEN_2064 & _GEN_2032) begin // @[cache.scala 84:50]
          tagArray_0_15 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_0 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1552) begin // @[cache.scala 84:50]
          tagArray_1_0 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_1 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1584) begin // @[cache.scala 84:50]
          tagArray_1_1 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_2 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1616) begin // @[cache.scala 84:50]
          tagArray_1_2 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_3 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1648) begin // @[cache.scala 84:50]
          tagArray_1_3 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_4 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1680) begin // @[cache.scala 84:50]
          tagArray_1_4 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_5 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1712) begin // @[cache.scala 84:50]
          tagArray_1_5 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_6 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1744) begin // @[cache.scala 84:50]
          tagArray_1_6 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_7 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1776) begin // @[cache.scala 84:50]
          tagArray_1_7 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_8 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1808) begin // @[cache.scala 84:50]
          tagArray_1_8 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_9 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1840) begin // @[cache.scala 84:50]
          tagArray_1_9 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_10 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1872) begin // @[cache.scala 84:50]
          tagArray_1_10 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_11 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1904) begin // @[cache.scala 84:50]
          tagArray_1_11 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_12 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1936) begin // @[cache.scala 84:50]
          tagArray_1_12 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_13 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_1968) begin // @[cache.scala 84:50]
          tagArray_1_13 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_14 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_2000) begin // @[cache.scala 84:50]
          tagArray_1_14 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 31:29]
      tagArray_1_15 <= 22'h0; // @[cache.scala 31:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        if (replace_set & _GEN_2032) begin // @[cache.scala 84:50]
          tagArray_1_15 <= tag; // @[cache.scala 84:50]
        end
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_0 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_0 <= _GEN_589;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_1 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_1 <= _GEN_590;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_2 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_2 <= _GEN_591;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_3 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_3 <= _GEN_592;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_4 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_4 <= _GEN_593;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_5 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_5 <= _GEN_594;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_6 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_6 <= _GEN_595;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_7 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_7 <= _GEN_596;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_8 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_8 <= _GEN_597;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_9 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_9 <= _GEN_598;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_10 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_10 <= _GEN_599;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_11 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_11 <= _GEN_600;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_12 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_12 <= _GEN_601;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_13 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_13 <= _GEN_602;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_14 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_14 <= _GEN_603;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_0_15 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_0_15 <= _GEN_604;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_0 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_0 <= _GEN_605;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_1 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_1 <= _GEN_606;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_2 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_2 <= _GEN_607;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_3 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_3 <= _GEN_608;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_4 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_4 <= _GEN_609;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_5 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_5 <= _GEN_610;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_6 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_6 <= _GEN_611;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_7 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_7 <= _GEN_612;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_8 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_8 <= _GEN_613;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_9 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_9 <= _GEN_614;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_10 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_10 <= _GEN_615;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_11 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_11 <= _GEN_616;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_12 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_12 <= _GEN_617;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_13 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_13 <= _GEN_618;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_14 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_14 <= _GEN_619;
      end
    end
    if (reset) begin // @[cache.scala 32:29]
      validArray_1_15 <= 1'h0; // @[cache.scala 32:29]
    end else if (state_cache == 3'h3 & _off_T) begin // @[cache.scala 80:58]
      if (to_sram_r_bits_last) begin // @[cache.scala 82:35]
        validArray_1_15 <= _GEN_620;
      end
    end
    if (reset) begin // @[cache.scala 45:24]
      off <= 4'h0; // @[cache.scala 45:24]
    end else if (!(3'h0 == state_cache)) begin // @[cache.scala 49:26]
      if (!(3'h1 == state_cache)) begin // @[cache.scala 49:26]
        if (3'h2 == state_cache) begin // @[cache.scala 49:26]
          off <= 4'h0; // @[cache.scala 63:25]
        end else begin
          off <= _GEN_67;
        end
      end
    end
    if (reset) begin // @[cache.scala 48:30]
      state_cache <= 3'h0; // @[cache.scala 48:30]
    end else if (3'h0 == state_cache) begin // @[cache.scala 49:26]
      if (_T_1) begin // @[cache.scala 51:34]
        if (hit) begin // @[cache.scala 52:35]
          state_cache <= 3'h1;
        end else begin
          state_cache <= 3'h2;
        end
      end else begin
        state_cache <= 3'h0; // @[cache.scala 54:29]
      end
    end else if (3'h1 == state_cache) begin // @[cache.scala 49:26]
      state_cache <= 3'h0; // @[cache.scala 58:25]
    end else if (3'h2 == state_cache) begin // @[cache.scala 49:26]
      state_cache <= _state_cache_T_2; // @[cache.scala 62:25]
    end else begin
      state_cache <= _GEN_66;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_0[initvar] = _RAND_0[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_1[initvar] = _RAND_3[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_2[initvar] = _RAND_6[31:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_3[initvar] = _RAND_9[31:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_4[initvar] = _RAND_12[31:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_5[initvar] = _RAND_15[31:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_6[initvar] = _RAND_18[31:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_7[initvar] = _RAND_21[31:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_8[initvar] = _RAND_24[31:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_9[initvar] = _RAND_27[31:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_10[initvar] = _RAND_30[31:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_11[initvar] = _RAND_33[31:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_12[initvar] = _RAND_36[31:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_13[initvar] = _RAND_39[31:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_14[initvar] = _RAND_42[31:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_0_15[initvar] = _RAND_45[31:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_0[initvar] = _RAND_48[31:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_1[initvar] = _RAND_51[31:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_2[initvar] = _RAND_54[31:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_3[initvar] = _RAND_57[31:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_4[initvar] = _RAND_60[31:0];
  _RAND_63 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_5[initvar] = _RAND_63[31:0];
  _RAND_66 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_6[initvar] = _RAND_66[31:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_7[initvar] = _RAND_69[31:0];
  _RAND_72 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_8[initvar] = _RAND_72[31:0];
  _RAND_75 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_9[initvar] = _RAND_75[31:0];
  _RAND_78 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_10[initvar] = _RAND_78[31:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_11[initvar] = _RAND_81[31:0];
  _RAND_84 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_12[initvar] = _RAND_84[31:0];
  _RAND_87 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_13[initvar] = _RAND_87[31:0];
  _RAND_90 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_14[initvar] = _RAND_90[31:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_1_15[initvar] = _RAND_93[31:0];
  _RAND_96 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_0[initvar] = _RAND_96[31:0];
  _RAND_99 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_1[initvar] = _RAND_99[31:0];
  _RAND_102 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_2[initvar] = _RAND_102[31:0];
  _RAND_105 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_3[initvar] = _RAND_105[31:0];
  _RAND_108 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_4[initvar] = _RAND_108[31:0];
  _RAND_111 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_5[initvar] = _RAND_111[31:0];
  _RAND_114 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_6[initvar] = _RAND_114[31:0];
  _RAND_117 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_7[initvar] = _RAND_117[31:0];
  _RAND_120 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_8[initvar] = _RAND_120[31:0];
  _RAND_123 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_9[initvar] = _RAND_123[31:0];
  _RAND_126 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_10[initvar] = _RAND_126[31:0];
  _RAND_129 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_11[initvar] = _RAND_129[31:0];
  _RAND_132 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_12[initvar] = _RAND_132[31:0];
  _RAND_135 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_13[initvar] = _RAND_135[31:0];
  _RAND_138 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_14[initvar] = _RAND_138[31:0];
  _RAND_141 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_2_15[initvar] = _RAND_141[31:0];
  _RAND_144 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_0[initvar] = _RAND_144[31:0];
  _RAND_147 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_1[initvar] = _RAND_147[31:0];
  _RAND_150 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_2[initvar] = _RAND_150[31:0];
  _RAND_153 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_3[initvar] = _RAND_153[31:0];
  _RAND_156 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_4[initvar] = _RAND_156[31:0];
  _RAND_159 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_5[initvar] = _RAND_159[31:0];
  _RAND_162 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_6[initvar] = _RAND_162[31:0];
  _RAND_165 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_7[initvar] = _RAND_165[31:0];
  _RAND_168 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_8[initvar] = _RAND_168[31:0];
  _RAND_171 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_9[initvar] = _RAND_171[31:0];
  _RAND_174 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_10[initvar] = _RAND_174[31:0];
  _RAND_177 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_11[initvar] = _RAND_177[31:0];
  _RAND_180 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_12[initvar] = _RAND_180[31:0];
  _RAND_183 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_13[initvar] = _RAND_183[31:0];
  _RAND_186 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_14[initvar] = _RAND_186[31:0];
  _RAND_189 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_3_15[initvar] = _RAND_189[31:0];
  _RAND_192 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_0[initvar] = _RAND_192[31:0];
  _RAND_195 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_1[initvar] = _RAND_195[31:0];
  _RAND_198 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_2[initvar] = _RAND_198[31:0];
  _RAND_201 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_3[initvar] = _RAND_201[31:0];
  _RAND_204 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_4[initvar] = _RAND_204[31:0];
  _RAND_207 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_5[initvar] = _RAND_207[31:0];
  _RAND_210 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_6[initvar] = _RAND_210[31:0];
  _RAND_213 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_7[initvar] = _RAND_213[31:0];
  _RAND_216 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_8[initvar] = _RAND_216[31:0];
  _RAND_219 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_9[initvar] = _RAND_219[31:0];
  _RAND_222 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_10[initvar] = _RAND_222[31:0];
  _RAND_225 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_11[initvar] = _RAND_225[31:0];
  _RAND_228 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_12[initvar] = _RAND_228[31:0];
  _RAND_231 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_13[initvar] = _RAND_231[31:0];
  _RAND_234 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_14[initvar] = _RAND_234[31:0];
  _RAND_237 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_4_15[initvar] = _RAND_237[31:0];
  _RAND_240 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_0[initvar] = _RAND_240[31:0];
  _RAND_243 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_1[initvar] = _RAND_243[31:0];
  _RAND_246 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_2[initvar] = _RAND_246[31:0];
  _RAND_249 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_3[initvar] = _RAND_249[31:0];
  _RAND_252 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_4[initvar] = _RAND_252[31:0];
  _RAND_255 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_5[initvar] = _RAND_255[31:0];
  _RAND_258 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_6[initvar] = _RAND_258[31:0];
  _RAND_261 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_7[initvar] = _RAND_261[31:0];
  _RAND_264 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_8[initvar] = _RAND_264[31:0];
  _RAND_267 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_9[initvar] = _RAND_267[31:0];
  _RAND_270 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_10[initvar] = _RAND_270[31:0];
  _RAND_273 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_11[initvar] = _RAND_273[31:0];
  _RAND_276 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_12[initvar] = _RAND_276[31:0];
  _RAND_279 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_13[initvar] = _RAND_279[31:0];
  _RAND_282 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_14[initvar] = _RAND_282[31:0];
  _RAND_285 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_5_15[initvar] = _RAND_285[31:0];
  _RAND_288 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_0[initvar] = _RAND_288[31:0];
  _RAND_291 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_1[initvar] = _RAND_291[31:0];
  _RAND_294 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_2[initvar] = _RAND_294[31:0];
  _RAND_297 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_3[initvar] = _RAND_297[31:0];
  _RAND_300 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_4[initvar] = _RAND_300[31:0];
  _RAND_303 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_5[initvar] = _RAND_303[31:0];
  _RAND_306 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_6[initvar] = _RAND_306[31:0];
  _RAND_309 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_7[initvar] = _RAND_309[31:0];
  _RAND_312 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_8[initvar] = _RAND_312[31:0];
  _RAND_315 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_9[initvar] = _RAND_315[31:0];
  _RAND_318 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_10[initvar] = _RAND_318[31:0];
  _RAND_321 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_11[initvar] = _RAND_321[31:0];
  _RAND_324 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_12[initvar] = _RAND_324[31:0];
  _RAND_327 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_13[initvar] = _RAND_327[31:0];
  _RAND_330 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_14[initvar] = _RAND_330[31:0];
  _RAND_333 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_6_15[initvar] = _RAND_333[31:0];
  _RAND_336 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_0[initvar] = _RAND_336[31:0];
  _RAND_339 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_1[initvar] = _RAND_339[31:0];
  _RAND_342 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_2[initvar] = _RAND_342[31:0];
  _RAND_345 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_3[initvar] = _RAND_345[31:0];
  _RAND_348 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_4[initvar] = _RAND_348[31:0];
  _RAND_351 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_5[initvar] = _RAND_351[31:0];
  _RAND_354 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_6[initvar] = _RAND_354[31:0];
  _RAND_357 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_7[initvar] = _RAND_357[31:0];
  _RAND_360 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_8[initvar] = _RAND_360[31:0];
  _RAND_363 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_9[initvar] = _RAND_363[31:0];
  _RAND_366 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_10[initvar] = _RAND_366[31:0];
  _RAND_369 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_11[initvar] = _RAND_369[31:0];
  _RAND_372 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_12[initvar] = _RAND_372[31:0];
  _RAND_375 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_13[initvar] = _RAND_375[31:0];
  _RAND_378 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_14[initvar] = _RAND_378[31:0];
  _RAND_381 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_7_15[initvar] = _RAND_381[31:0];
  _RAND_384 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_0[initvar] = _RAND_384[31:0];
  _RAND_387 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_1[initvar] = _RAND_387[31:0];
  _RAND_390 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_2[initvar] = _RAND_390[31:0];
  _RAND_393 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_3[initvar] = _RAND_393[31:0];
  _RAND_396 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_4[initvar] = _RAND_396[31:0];
  _RAND_399 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_5[initvar] = _RAND_399[31:0];
  _RAND_402 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_6[initvar] = _RAND_402[31:0];
  _RAND_405 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_7[initvar] = _RAND_405[31:0];
  _RAND_408 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_8[initvar] = _RAND_408[31:0];
  _RAND_411 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_9[initvar] = _RAND_411[31:0];
  _RAND_414 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_10[initvar] = _RAND_414[31:0];
  _RAND_417 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_11[initvar] = _RAND_417[31:0];
  _RAND_420 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_12[initvar] = _RAND_420[31:0];
  _RAND_423 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_13[initvar] = _RAND_423[31:0];
  _RAND_426 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_14[initvar] = _RAND_426[31:0];
  _RAND_429 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_8_15[initvar] = _RAND_429[31:0];
  _RAND_432 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_0[initvar] = _RAND_432[31:0];
  _RAND_435 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_1[initvar] = _RAND_435[31:0];
  _RAND_438 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_2[initvar] = _RAND_438[31:0];
  _RAND_441 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_3[initvar] = _RAND_441[31:0];
  _RAND_444 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_4[initvar] = _RAND_444[31:0];
  _RAND_447 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_5[initvar] = _RAND_447[31:0];
  _RAND_450 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_6[initvar] = _RAND_450[31:0];
  _RAND_453 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_7[initvar] = _RAND_453[31:0];
  _RAND_456 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_8[initvar] = _RAND_456[31:0];
  _RAND_459 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_9[initvar] = _RAND_459[31:0];
  _RAND_462 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_10[initvar] = _RAND_462[31:0];
  _RAND_465 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_11[initvar] = _RAND_465[31:0];
  _RAND_468 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_12[initvar] = _RAND_468[31:0];
  _RAND_471 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_13[initvar] = _RAND_471[31:0];
  _RAND_474 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_14[initvar] = _RAND_474[31:0];
  _RAND_477 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_9_15[initvar] = _RAND_477[31:0];
  _RAND_480 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_0[initvar] = _RAND_480[31:0];
  _RAND_483 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_1[initvar] = _RAND_483[31:0];
  _RAND_486 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_2[initvar] = _RAND_486[31:0];
  _RAND_489 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_3[initvar] = _RAND_489[31:0];
  _RAND_492 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_4[initvar] = _RAND_492[31:0];
  _RAND_495 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_5[initvar] = _RAND_495[31:0];
  _RAND_498 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_6[initvar] = _RAND_498[31:0];
  _RAND_501 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_7[initvar] = _RAND_501[31:0];
  _RAND_504 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_8[initvar] = _RAND_504[31:0];
  _RAND_507 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_9[initvar] = _RAND_507[31:0];
  _RAND_510 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_10[initvar] = _RAND_510[31:0];
  _RAND_513 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_11[initvar] = _RAND_513[31:0];
  _RAND_516 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_12[initvar] = _RAND_516[31:0];
  _RAND_519 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_13[initvar] = _RAND_519[31:0];
  _RAND_522 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_14[initvar] = _RAND_522[31:0];
  _RAND_525 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_10_15[initvar] = _RAND_525[31:0];
  _RAND_528 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_0[initvar] = _RAND_528[31:0];
  _RAND_531 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_1[initvar] = _RAND_531[31:0];
  _RAND_534 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_2[initvar] = _RAND_534[31:0];
  _RAND_537 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_3[initvar] = _RAND_537[31:0];
  _RAND_540 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_4[initvar] = _RAND_540[31:0];
  _RAND_543 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_5[initvar] = _RAND_543[31:0];
  _RAND_546 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_6[initvar] = _RAND_546[31:0];
  _RAND_549 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_7[initvar] = _RAND_549[31:0];
  _RAND_552 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_8[initvar] = _RAND_552[31:0];
  _RAND_555 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_9[initvar] = _RAND_555[31:0];
  _RAND_558 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_10[initvar] = _RAND_558[31:0];
  _RAND_561 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_11[initvar] = _RAND_561[31:0];
  _RAND_564 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_12[initvar] = _RAND_564[31:0];
  _RAND_567 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_13[initvar] = _RAND_567[31:0];
  _RAND_570 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_14[initvar] = _RAND_570[31:0];
  _RAND_573 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_11_15[initvar] = _RAND_573[31:0];
  _RAND_576 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_0[initvar] = _RAND_576[31:0];
  _RAND_579 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_1[initvar] = _RAND_579[31:0];
  _RAND_582 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_2[initvar] = _RAND_582[31:0];
  _RAND_585 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_3[initvar] = _RAND_585[31:0];
  _RAND_588 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_4[initvar] = _RAND_588[31:0];
  _RAND_591 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_5[initvar] = _RAND_591[31:0];
  _RAND_594 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_6[initvar] = _RAND_594[31:0];
  _RAND_597 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_7[initvar] = _RAND_597[31:0];
  _RAND_600 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_8[initvar] = _RAND_600[31:0];
  _RAND_603 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_9[initvar] = _RAND_603[31:0];
  _RAND_606 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_10[initvar] = _RAND_606[31:0];
  _RAND_609 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_11[initvar] = _RAND_609[31:0];
  _RAND_612 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_12[initvar] = _RAND_612[31:0];
  _RAND_615 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_13[initvar] = _RAND_615[31:0];
  _RAND_618 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_14[initvar] = _RAND_618[31:0];
  _RAND_621 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_12_15[initvar] = _RAND_621[31:0];
  _RAND_624 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_0[initvar] = _RAND_624[31:0];
  _RAND_627 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_1[initvar] = _RAND_627[31:0];
  _RAND_630 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_2[initvar] = _RAND_630[31:0];
  _RAND_633 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_3[initvar] = _RAND_633[31:0];
  _RAND_636 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_4[initvar] = _RAND_636[31:0];
  _RAND_639 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_5[initvar] = _RAND_639[31:0];
  _RAND_642 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_6[initvar] = _RAND_642[31:0];
  _RAND_645 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_7[initvar] = _RAND_645[31:0];
  _RAND_648 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_8[initvar] = _RAND_648[31:0];
  _RAND_651 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_9[initvar] = _RAND_651[31:0];
  _RAND_654 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_10[initvar] = _RAND_654[31:0];
  _RAND_657 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_11[initvar] = _RAND_657[31:0];
  _RAND_660 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_12[initvar] = _RAND_660[31:0];
  _RAND_663 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_13[initvar] = _RAND_663[31:0];
  _RAND_666 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_14[initvar] = _RAND_666[31:0];
  _RAND_669 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_13_15[initvar] = _RAND_669[31:0];
  _RAND_672 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_0[initvar] = _RAND_672[31:0];
  _RAND_675 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_1[initvar] = _RAND_675[31:0];
  _RAND_678 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_2[initvar] = _RAND_678[31:0];
  _RAND_681 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_3[initvar] = _RAND_681[31:0];
  _RAND_684 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_4[initvar] = _RAND_684[31:0];
  _RAND_687 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_5[initvar] = _RAND_687[31:0];
  _RAND_690 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_6[initvar] = _RAND_690[31:0];
  _RAND_693 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_7[initvar] = _RAND_693[31:0];
  _RAND_696 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_8[initvar] = _RAND_696[31:0];
  _RAND_699 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_9[initvar] = _RAND_699[31:0];
  _RAND_702 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_10[initvar] = _RAND_702[31:0];
  _RAND_705 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_11[initvar] = _RAND_705[31:0];
  _RAND_708 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_12[initvar] = _RAND_708[31:0];
  _RAND_711 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_13[initvar] = _RAND_711[31:0];
  _RAND_714 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_14[initvar] = _RAND_714[31:0];
  _RAND_717 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_14_15[initvar] = _RAND_717[31:0];
  _RAND_720 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_0[initvar] = _RAND_720[31:0];
  _RAND_723 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_1[initvar] = _RAND_723[31:0];
  _RAND_726 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_2[initvar] = _RAND_726[31:0];
  _RAND_729 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_3[initvar] = _RAND_729[31:0];
  _RAND_732 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_4[initvar] = _RAND_732[31:0];
  _RAND_735 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_5[initvar] = _RAND_735[31:0];
  _RAND_738 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_6[initvar] = _RAND_738[31:0];
  _RAND_741 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_7[initvar] = _RAND_741[31:0];
  _RAND_744 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_8[initvar] = _RAND_744[31:0];
  _RAND_747 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_9[initvar] = _RAND_747[31:0];
  _RAND_750 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_10[initvar] = _RAND_750[31:0];
  _RAND_753 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_11[initvar] = _RAND_753[31:0];
  _RAND_756 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_12[initvar] = _RAND_756[31:0];
  _RAND_759 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_13[initvar] = _RAND_759[31:0];
  _RAND_762 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_14[initvar] = _RAND_762[31:0];
  _RAND_765 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataArray_15_15[initvar] = _RAND_765[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  dataArray_0_0_cachedata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  dataArray_0_0_cachedata_MPORT_addr_pipe_0 = _RAND_2[0:0];
  _RAND_4 = {1{`RANDOM}};
  dataArray_0_1_cachedata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataArray_0_1_cachedata_MPORT_addr_pipe_0 = _RAND_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataArray_0_2_cachedata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataArray_0_2_cachedata_MPORT_addr_pipe_0 = _RAND_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  dataArray_0_3_cachedata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataArray_0_3_cachedata_MPORT_addr_pipe_0 = _RAND_11[0:0];
  _RAND_13 = {1{`RANDOM}};
  dataArray_0_4_cachedata_MPORT_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataArray_0_4_cachedata_MPORT_addr_pipe_0 = _RAND_14[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataArray_0_5_cachedata_MPORT_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dataArray_0_5_cachedata_MPORT_addr_pipe_0 = _RAND_17[0:0];
  _RAND_19 = {1{`RANDOM}};
  dataArray_0_6_cachedata_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dataArray_0_6_cachedata_MPORT_addr_pipe_0 = _RAND_20[0:0];
  _RAND_22 = {1{`RANDOM}};
  dataArray_0_7_cachedata_MPORT_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  dataArray_0_7_cachedata_MPORT_addr_pipe_0 = _RAND_23[0:0];
  _RAND_25 = {1{`RANDOM}};
  dataArray_0_8_cachedata_MPORT_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  dataArray_0_8_cachedata_MPORT_addr_pipe_0 = _RAND_26[0:0];
  _RAND_28 = {1{`RANDOM}};
  dataArray_0_9_cachedata_MPORT_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dataArray_0_9_cachedata_MPORT_addr_pipe_0 = _RAND_29[0:0];
  _RAND_31 = {1{`RANDOM}};
  dataArray_0_10_cachedata_MPORT_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataArray_0_10_cachedata_MPORT_addr_pipe_0 = _RAND_32[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataArray_0_11_cachedata_MPORT_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataArray_0_11_cachedata_MPORT_addr_pipe_0 = _RAND_35[0:0];
  _RAND_37 = {1{`RANDOM}};
  dataArray_0_12_cachedata_MPORT_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataArray_0_12_cachedata_MPORT_addr_pipe_0 = _RAND_38[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataArray_0_13_cachedata_MPORT_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dataArray_0_13_cachedata_MPORT_addr_pipe_0 = _RAND_41[0:0];
  _RAND_43 = {1{`RANDOM}};
  dataArray_0_14_cachedata_MPORT_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dataArray_0_14_cachedata_MPORT_addr_pipe_0 = _RAND_44[0:0];
  _RAND_46 = {1{`RANDOM}};
  dataArray_0_15_cachedata_MPORT_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dataArray_0_15_cachedata_MPORT_addr_pipe_0 = _RAND_47[0:0];
  _RAND_49 = {1{`RANDOM}};
  dataArray_1_0_cachedata_MPORT_en_pipe_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dataArray_1_0_cachedata_MPORT_addr_pipe_0 = _RAND_50[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataArray_1_1_cachedata_MPORT_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dataArray_1_1_cachedata_MPORT_addr_pipe_0 = _RAND_53[0:0];
  _RAND_55 = {1{`RANDOM}};
  dataArray_1_2_cachedata_MPORT_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dataArray_1_2_cachedata_MPORT_addr_pipe_0 = _RAND_56[0:0];
  _RAND_58 = {1{`RANDOM}};
  dataArray_1_3_cachedata_MPORT_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dataArray_1_3_cachedata_MPORT_addr_pipe_0 = _RAND_59[0:0];
  _RAND_61 = {1{`RANDOM}};
  dataArray_1_4_cachedata_MPORT_en_pipe_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dataArray_1_4_cachedata_MPORT_addr_pipe_0 = _RAND_62[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataArray_1_5_cachedata_MPORT_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dataArray_1_5_cachedata_MPORT_addr_pipe_0 = _RAND_65[0:0];
  _RAND_67 = {1{`RANDOM}};
  dataArray_1_6_cachedata_MPORT_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dataArray_1_6_cachedata_MPORT_addr_pipe_0 = _RAND_68[0:0];
  _RAND_70 = {1{`RANDOM}};
  dataArray_1_7_cachedata_MPORT_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dataArray_1_7_cachedata_MPORT_addr_pipe_0 = _RAND_71[0:0];
  _RAND_73 = {1{`RANDOM}};
  dataArray_1_8_cachedata_MPORT_en_pipe_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dataArray_1_8_cachedata_MPORT_addr_pipe_0 = _RAND_74[0:0];
  _RAND_76 = {1{`RANDOM}};
  dataArray_1_9_cachedata_MPORT_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dataArray_1_9_cachedata_MPORT_addr_pipe_0 = _RAND_77[0:0];
  _RAND_79 = {1{`RANDOM}};
  dataArray_1_10_cachedata_MPORT_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataArray_1_10_cachedata_MPORT_addr_pipe_0 = _RAND_80[0:0];
  _RAND_82 = {1{`RANDOM}};
  dataArray_1_11_cachedata_MPORT_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dataArray_1_11_cachedata_MPORT_addr_pipe_0 = _RAND_83[0:0];
  _RAND_85 = {1{`RANDOM}};
  dataArray_1_12_cachedata_MPORT_en_pipe_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dataArray_1_12_cachedata_MPORT_addr_pipe_0 = _RAND_86[0:0];
  _RAND_88 = {1{`RANDOM}};
  dataArray_1_13_cachedata_MPORT_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dataArray_1_13_cachedata_MPORT_addr_pipe_0 = _RAND_89[0:0];
  _RAND_91 = {1{`RANDOM}};
  dataArray_1_14_cachedata_MPORT_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dataArray_1_14_cachedata_MPORT_addr_pipe_0 = _RAND_92[0:0];
  _RAND_94 = {1{`RANDOM}};
  dataArray_1_15_cachedata_MPORT_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dataArray_1_15_cachedata_MPORT_addr_pipe_0 = _RAND_95[0:0];
  _RAND_97 = {1{`RANDOM}};
  dataArray_2_0_cachedata_MPORT_en_pipe_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dataArray_2_0_cachedata_MPORT_addr_pipe_0 = _RAND_98[0:0];
  _RAND_100 = {1{`RANDOM}};
  dataArray_2_1_cachedata_MPORT_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dataArray_2_1_cachedata_MPORT_addr_pipe_0 = _RAND_101[0:0];
  _RAND_103 = {1{`RANDOM}};
  dataArray_2_2_cachedata_MPORT_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dataArray_2_2_cachedata_MPORT_addr_pipe_0 = _RAND_104[0:0];
  _RAND_106 = {1{`RANDOM}};
  dataArray_2_3_cachedata_MPORT_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dataArray_2_3_cachedata_MPORT_addr_pipe_0 = _RAND_107[0:0];
  _RAND_109 = {1{`RANDOM}};
  dataArray_2_4_cachedata_MPORT_en_pipe_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dataArray_2_4_cachedata_MPORT_addr_pipe_0 = _RAND_110[0:0];
  _RAND_112 = {1{`RANDOM}};
  dataArray_2_5_cachedata_MPORT_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dataArray_2_5_cachedata_MPORT_addr_pipe_0 = _RAND_113[0:0];
  _RAND_115 = {1{`RANDOM}};
  dataArray_2_6_cachedata_MPORT_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dataArray_2_6_cachedata_MPORT_addr_pipe_0 = _RAND_116[0:0];
  _RAND_118 = {1{`RANDOM}};
  dataArray_2_7_cachedata_MPORT_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dataArray_2_7_cachedata_MPORT_addr_pipe_0 = _RAND_119[0:0];
  _RAND_121 = {1{`RANDOM}};
  dataArray_2_8_cachedata_MPORT_en_pipe_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dataArray_2_8_cachedata_MPORT_addr_pipe_0 = _RAND_122[0:0];
  _RAND_124 = {1{`RANDOM}};
  dataArray_2_9_cachedata_MPORT_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dataArray_2_9_cachedata_MPORT_addr_pipe_0 = _RAND_125[0:0];
  _RAND_127 = {1{`RANDOM}};
  dataArray_2_10_cachedata_MPORT_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dataArray_2_10_cachedata_MPORT_addr_pipe_0 = _RAND_128[0:0];
  _RAND_130 = {1{`RANDOM}};
  dataArray_2_11_cachedata_MPORT_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  dataArray_2_11_cachedata_MPORT_addr_pipe_0 = _RAND_131[0:0];
  _RAND_133 = {1{`RANDOM}};
  dataArray_2_12_cachedata_MPORT_en_pipe_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  dataArray_2_12_cachedata_MPORT_addr_pipe_0 = _RAND_134[0:0];
  _RAND_136 = {1{`RANDOM}};
  dataArray_2_13_cachedata_MPORT_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dataArray_2_13_cachedata_MPORT_addr_pipe_0 = _RAND_137[0:0];
  _RAND_139 = {1{`RANDOM}};
  dataArray_2_14_cachedata_MPORT_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dataArray_2_14_cachedata_MPORT_addr_pipe_0 = _RAND_140[0:0];
  _RAND_142 = {1{`RANDOM}};
  dataArray_2_15_cachedata_MPORT_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dataArray_2_15_cachedata_MPORT_addr_pipe_0 = _RAND_143[0:0];
  _RAND_145 = {1{`RANDOM}};
  dataArray_3_0_cachedata_MPORT_en_pipe_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dataArray_3_0_cachedata_MPORT_addr_pipe_0 = _RAND_146[0:0];
  _RAND_148 = {1{`RANDOM}};
  dataArray_3_1_cachedata_MPORT_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dataArray_3_1_cachedata_MPORT_addr_pipe_0 = _RAND_149[0:0];
  _RAND_151 = {1{`RANDOM}};
  dataArray_3_2_cachedata_MPORT_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dataArray_3_2_cachedata_MPORT_addr_pipe_0 = _RAND_152[0:0];
  _RAND_154 = {1{`RANDOM}};
  dataArray_3_3_cachedata_MPORT_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dataArray_3_3_cachedata_MPORT_addr_pipe_0 = _RAND_155[0:0];
  _RAND_157 = {1{`RANDOM}};
  dataArray_3_4_cachedata_MPORT_en_pipe_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dataArray_3_4_cachedata_MPORT_addr_pipe_0 = _RAND_158[0:0];
  _RAND_160 = {1{`RANDOM}};
  dataArray_3_5_cachedata_MPORT_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dataArray_3_5_cachedata_MPORT_addr_pipe_0 = _RAND_161[0:0];
  _RAND_163 = {1{`RANDOM}};
  dataArray_3_6_cachedata_MPORT_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dataArray_3_6_cachedata_MPORT_addr_pipe_0 = _RAND_164[0:0];
  _RAND_166 = {1{`RANDOM}};
  dataArray_3_7_cachedata_MPORT_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dataArray_3_7_cachedata_MPORT_addr_pipe_0 = _RAND_167[0:0];
  _RAND_169 = {1{`RANDOM}};
  dataArray_3_8_cachedata_MPORT_en_pipe_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dataArray_3_8_cachedata_MPORT_addr_pipe_0 = _RAND_170[0:0];
  _RAND_172 = {1{`RANDOM}};
  dataArray_3_9_cachedata_MPORT_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dataArray_3_9_cachedata_MPORT_addr_pipe_0 = _RAND_173[0:0];
  _RAND_175 = {1{`RANDOM}};
  dataArray_3_10_cachedata_MPORT_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dataArray_3_10_cachedata_MPORT_addr_pipe_0 = _RAND_176[0:0];
  _RAND_178 = {1{`RANDOM}};
  dataArray_3_11_cachedata_MPORT_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dataArray_3_11_cachedata_MPORT_addr_pipe_0 = _RAND_179[0:0];
  _RAND_181 = {1{`RANDOM}};
  dataArray_3_12_cachedata_MPORT_en_pipe_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dataArray_3_12_cachedata_MPORT_addr_pipe_0 = _RAND_182[0:0];
  _RAND_184 = {1{`RANDOM}};
  dataArray_3_13_cachedata_MPORT_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dataArray_3_13_cachedata_MPORT_addr_pipe_0 = _RAND_185[0:0];
  _RAND_187 = {1{`RANDOM}};
  dataArray_3_14_cachedata_MPORT_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dataArray_3_14_cachedata_MPORT_addr_pipe_0 = _RAND_188[0:0];
  _RAND_190 = {1{`RANDOM}};
  dataArray_3_15_cachedata_MPORT_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dataArray_3_15_cachedata_MPORT_addr_pipe_0 = _RAND_191[0:0];
  _RAND_193 = {1{`RANDOM}};
  dataArray_4_0_cachedata_MPORT_en_pipe_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dataArray_4_0_cachedata_MPORT_addr_pipe_0 = _RAND_194[0:0];
  _RAND_196 = {1{`RANDOM}};
  dataArray_4_1_cachedata_MPORT_en_pipe_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dataArray_4_1_cachedata_MPORT_addr_pipe_0 = _RAND_197[0:0];
  _RAND_199 = {1{`RANDOM}};
  dataArray_4_2_cachedata_MPORT_en_pipe_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dataArray_4_2_cachedata_MPORT_addr_pipe_0 = _RAND_200[0:0];
  _RAND_202 = {1{`RANDOM}};
  dataArray_4_3_cachedata_MPORT_en_pipe_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dataArray_4_3_cachedata_MPORT_addr_pipe_0 = _RAND_203[0:0];
  _RAND_205 = {1{`RANDOM}};
  dataArray_4_4_cachedata_MPORT_en_pipe_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dataArray_4_4_cachedata_MPORT_addr_pipe_0 = _RAND_206[0:0];
  _RAND_208 = {1{`RANDOM}};
  dataArray_4_5_cachedata_MPORT_en_pipe_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dataArray_4_5_cachedata_MPORT_addr_pipe_0 = _RAND_209[0:0];
  _RAND_211 = {1{`RANDOM}};
  dataArray_4_6_cachedata_MPORT_en_pipe_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dataArray_4_6_cachedata_MPORT_addr_pipe_0 = _RAND_212[0:0];
  _RAND_214 = {1{`RANDOM}};
  dataArray_4_7_cachedata_MPORT_en_pipe_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dataArray_4_7_cachedata_MPORT_addr_pipe_0 = _RAND_215[0:0];
  _RAND_217 = {1{`RANDOM}};
  dataArray_4_8_cachedata_MPORT_en_pipe_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dataArray_4_8_cachedata_MPORT_addr_pipe_0 = _RAND_218[0:0];
  _RAND_220 = {1{`RANDOM}};
  dataArray_4_9_cachedata_MPORT_en_pipe_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dataArray_4_9_cachedata_MPORT_addr_pipe_0 = _RAND_221[0:0];
  _RAND_223 = {1{`RANDOM}};
  dataArray_4_10_cachedata_MPORT_en_pipe_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dataArray_4_10_cachedata_MPORT_addr_pipe_0 = _RAND_224[0:0];
  _RAND_226 = {1{`RANDOM}};
  dataArray_4_11_cachedata_MPORT_en_pipe_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dataArray_4_11_cachedata_MPORT_addr_pipe_0 = _RAND_227[0:0];
  _RAND_229 = {1{`RANDOM}};
  dataArray_4_12_cachedata_MPORT_en_pipe_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dataArray_4_12_cachedata_MPORT_addr_pipe_0 = _RAND_230[0:0];
  _RAND_232 = {1{`RANDOM}};
  dataArray_4_13_cachedata_MPORT_en_pipe_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dataArray_4_13_cachedata_MPORT_addr_pipe_0 = _RAND_233[0:0];
  _RAND_235 = {1{`RANDOM}};
  dataArray_4_14_cachedata_MPORT_en_pipe_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dataArray_4_14_cachedata_MPORT_addr_pipe_0 = _RAND_236[0:0];
  _RAND_238 = {1{`RANDOM}};
  dataArray_4_15_cachedata_MPORT_en_pipe_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dataArray_4_15_cachedata_MPORT_addr_pipe_0 = _RAND_239[0:0];
  _RAND_241 = {1{`RANDOM}};
  dataArray_5_0_cachedata_MPORT_en_pipe_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dataArray_5_0_cachedata_MPORT_addr_pipe_0 = _RAND_242[0:0];
  _RAND_244 = {1{`RANDOM}};
  dataArray_5_1_cachedata_MPORT_en_pipe_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dataArray_5_1_cachedata_MPORT_addr_pipe_0 = _RAND_245[0:0];
  _RAND_247 = {1{`RANDOM}};
  dataArray_5_2_cachedata_MPORT_en_pipe_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dataArray_5_2_cachedata_MPORT_addr_pipe_0 = _RAND_248[0:0];
  _RAND_250 = {1{`RANDOM}};
  dataArray_5_3_cachedata_MPORT_en_pipe_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dataArray_5_3_cachedata_MPORT_addr_pipe_0 = _RAND_251[0:0];
  _RAND_253 = {1{`RANDOM}};
  dataArray_5_4_cachedata_MPORT_en_pipe_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dataArray_5_4_cachedata_MPORT_addr_pipe_0 = _RAND_254[0:0];
  _RAND_256 = {1{`RANDOM}};
  dataArray_5_5_cachedata_MPORT_en_pipe_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  dataArray_5_5_cachedata_MPORT_addr_pipe_0 = _RAND_257[0:0];
  _RAND_259 = {1{`RANDOM}};
  dataArray_5_6_cachedata_MPORT_en_pipe_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dataArray_5_6_cachedata_MPORT_addr_pipe_0 = _RAND_260[0:0];
  _RAND_262 = {1{`RANDOM}};
  dataArray_5_7_cachedata_MPORT_en_pipe_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  dataArray_5_7_cachedata_MPORT_addr_pipe_0 = _RAND_263[0:0];
  _RAND_265 = {1{`RANDOM}};
  dataArray_5_8_cachedata_MPORT_en_pipe_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  dataArray_5_8_cachedata_MPORT_addr_pipe_0 = _RAND_266[0:0];
  _RAND_268 = {1{`RANDOM}};
  dataArray_5_9_cachedata_MPORT_en_pipe_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  dataArray_5_9_cachedata_MPORT_addr_pipe_0 = _RAND_269[0:0];
  _RAND_271 = {1{`RANDOM}};
  dataArray_5_10_cachedata_MPORT_en_pipe_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  dataArray_5_10_cachedata_MPORT_addr_pipe_0 = _RAND_272[0:0];
  _RAND_274 = {1{`RANDOM}};
  dataArray_5_11_cachedata_MPORT_en_pipe_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  dataArray_5_11_cachedata_MPORT_addr_pipe_0 = _RAND_275[0:0];
  _RAND_277 = {1{`RANDOM}};
  dataArray_5_12_cachedata_MPORT_en_pipe_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  dataArray_5_12_cachedata_MPORT_addr_pipe_0 = _RAND_278[0:0];
  _RAND_280 = {1{`RANDOM}};
  dataArray_5_13_cachedata_MPORT_en_pipe_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  dataArray_5_13_cachedata_MPORT_addr_pipe_0 = _RAND_281[0:0];
  _RAND_283 = {1{`RANDOM}};
  dataArray_5_14_cachedata_MPORT_en_pipe_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  dataArray_5_14_cachedata_MPORT_addr_pipe_0 = _RAND_284[0:0];
  _RAND_286 = {1{`RANDOM}};
  dataArray_5_15_cachedata_MPORT_en_pipe_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  dataArray_5_15_cachedata_MPORT_addr_pipe_0 = _RAND_287[0:0];
  _RAND_289 = {1{`RANDOM}};
  dataArray_6_0_cachedata_MPORT_en_pipe_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  dataArray_6_0_cachedata_MPORT_addr_pipe_0 = _RAND_290[0:0];
  _RAND_292 = {1{`RANDOM}};
  dataArray_6_1_cachedata_MPORT_en_pipe_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  dataArray_6_1_cachedata_MPORT_addr_pipe_0 = _RAND_293[0:0];
  _RAND_295 = {1{`RANDOM}};
  dataArray_6_2_cachedata_MPORT_en_pipe_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  dataArray_6_2_cachedata_MPORT_addr_pipe_0 = _RAND_296[0:0];
  _RAND_298 = {1{`RANDOM}};
  dataArray_6_3_cachedata_MPORT_en_pipe_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  dataArray_6_3_cachedata_MPORT_addr_pipe_0 = _RAND_299[0:0];
  _RAND_301 = {1{`RANDOM}};
  dataArray_6_4_cachedata_MPORT_en_pipe_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  dataArray_6_4_cachedata_MPORT_addr_pipe_0 = _RAND_302[0:0];
  _RAND_304 = {1{`RANDOM}};
  dataArray_6_5_cachedata_MPORT_en_pipe_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  dataArray_6_5_cachedata_MPORT_addr_pipe_0 = _RAND_305[0:0];
  _RAND_307 = {1{`RANDOM}};
  dataArray_6_6_cachedata_MPORT_en_pipe_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  dataArray_6_6_cachedata_MPORT_addr_pipe_0 = _RAND_308[0:0];
  _RAND_310 = {1{`RANDOM}};
  dataArray_6_7_cachedata_MPORT_en_pipe_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  dataArray_6_7_cachedata_MPORT_addr_pipe_0 = _RAND_311[0:0];
  _RAND_313 = {1{`RANDOM}};
  dataArray_6_8_cachedata_MPORT_en_pipe_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  dataArray_6_8_cachedata_MPORT_addr_pipe_0 = _RAND_314[0:0];
  _RAND_316 = {1{`RANDOM}};
  dataArray_6_9_cachedata_MPORT_en_pipe_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  dataArray_6_9_cachedata_MPORT_addr_pipe_0 = _RAND_317[0:0];
  _RAND_319 = {1{`RANDOM}};
  dataArray_6_10_cachedata_MPORT_en_pipe_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  dataArray_6_10_cachedata_MPORT_addr_pipe_0 = _RAND_320[0:0];
  _RAND_322 = {1{`RANDOM}};
  dataArray_6_11_cachedata_MPORT_en_pipe_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  dataArray_6_11_cachedata_MPORT_addr_pipe_0 = _RAND_323[0:0];
  _RAND_325 = {1{`RANDOM}};
  dataArray_6_12_cachedata_MPORT_en_pipe_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  dataArray_6_12_cachedata_MPORT_addr_pipe_0 = _RAND_326[0:0];
  _RAND_328 = {1{`RANDOM}};
  dataArray_6_13_cachedata_MPORT_en_pipe_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  dataArray_6_13_cachedata_MPORT_addr_pipe_0 = _RAND_329[0:0];
  _RAND_331 = {1{`RANDOM}};
  dataArray_6_14_cachedata_MPORT_en_pipe_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  dataArray_6_14_cachedata_MPORT_addr_pipe_0 = _RAND_332[0:0];
  _RAND_334 = {1{`RANDOM}};
  dataArray_6_15_cachedata_MPORT_en_pipe_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  dataArray_6_15_cachedata_MPORT_addr_pipe_0 = _RAND_335[0:0];
  _RAND_337 = {1{`RANDOM}};
  dataArray_7_0_cachedata_MPORT_en_pipe_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dataArray_7_0_cachedata_MPORT_addr_pipe_0 = _RAND_338[0:0];
  _RAND_340 = {1{`RANDOM}};
  dataArray_7_1_cachedata_MPORT_en_pipe_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  dataArray_7_1_cachedata_MPORT_addr_pipe_0 = _RAND_341[0:0];
  _RAND_343 = {1{`RANDOM}};
  dataArray_7_2_cachedata_MPORT_en_pipe_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  dataArray_7_2_cachedata_MPORT_addr_pipe_0 = _RAND_344[0:0];
  _RAND_346 = {1{`RANDOM}};
  dataArray_7_3_cachedata_MPORT_en_pipe_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  dataArray_7_3_cachedata_MPORT_addr_pipe_0 = _RAND_347[0:0];
  _RAND_349 = {1{`RANDOM}};
  dataArray_7_4_cachedata_MPORT_en_pipe_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  dataArray_7_4_cachedata_MPORT_addr_pipe_0 = _RAND_350[0:0];
  _RAND_352 = {1{`RANDOM}};
  dataArray_7_5_cachedata_MPORT_en_pipe_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  dataArray_7_5_cachedata_MPORT_addr_pipe_0 = _RAND_353[0:0];
  _RAND_355 = {1{`RANDOM}};
  dataArray_7_6_cachedata_MPORT_en_pipe_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  dataArray_7_6_cachedata_MPORT_addr_pipe_0 = _RAND_356[0:0];
  _RAND_358 = {1{`RANDOM}};
  dataArray_7_7_cachedata_MPORT_en_pipe_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  dataArray_7_7_cachedata_MPORT_addr_pipe_0 = _RAND_359[0:0];
  _RAND_361 = {1{`RANDOM}};
  dataArray_7_8_cachedata_MPORT_en_pipe_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  dataArray_7_8_cachedata_MPORT_addr_pipe_0 = _RAND_362[0:0];
  _RAND_364 = {1{`RANDOM}};
  dataArray_7_9_cachedata_MPORT_en_pipe_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  dataArray_7_9_cachedata_MPORT_addr_pipe_0 = _RAND_365[0:0];
  _RAND_367 = {1{`RANDOM}};
  dataArray_7_10_cachedata_MPORT_en_pipe_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  dataArray_7_10_cachedata_MPORT_addr_pipe_0 = _RAND_368[0:0];
  _RAND_370 = {1{`RANDOM}};
  dataArray_7_11_cachedata_MPORT_en_pipe_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  dataArray_7_11_cachedata_MPORT_addr_pipe_0 = _RAND_371[0:0];
  _RAND_373 = {1{`RANDOM}};
  dataArray_7_12_cachedata_MPORT_en_pipe_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  dataArray_7_12_cachedata_MPORT_addr_pipe_0 = _RAND_374[0:0];
  _RAND_376 = {1{`RANDOM}};
  dataArray_7_13_cachedata_MPORT_en_pipe_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  dataArray_7_13_cachedata_MPORT_addr_pipe_0 = _RAND_377[0:0];
  _RAND_379 = {1{`RANDOM}};
  dataArray_7_14_cachedata_MPORT_en_pipe_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  dataArray_7_14_cachedata_MPORT_addr_pipe_0 = _RAND_380[0:0];
  _RAND_382 = {1{`RANDOM}};
  dataArray_7_15_cachedata_MPORT_en_pipe_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  dataArray_7_15_cachedata_MPORT_addr_pipe_0 = _RAND_383[0:0];
  _RAND_385 = {1{`RANDOM}};
  dataArray_8_0_cachedata_MPORT_en_pipe_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dataArray_8_0_cachedata_MPORT_addr_pipe_0 = _RAND_386[0:0];
  _RAND_388 = {1{`RANDOM}};
  dataArray_8_1_cachedata_MPORT_en_pipe_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dataArray_8_1_cachedata_MPORT_addr_pipe_0 = _RAND_389[0:0];
  _RAND_391 = {1{`RANDOM}};
  dataArray_8_2_cachedata_MPORT_en_pipe_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dataArray_8_2_cachedata_MPORT_addr_pipe_0 = _RAND_392[0:0];
  _RAND_394 = {1{`RANDOM}};
  dataArray_8_3_cachedata_MPORT_en_pipe_0 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dataArray_8_3_cachedata_MPORT_addr_pipe_0 = _RAND_395[0:0];
  _RAND_397 = {1{`RANDOM}};
  dataArray_8_4_cachedata_MPORT_en_pipe_0 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dataArray_8_4_cachedata_MPORT_addr_pipe_0 = _RAND_398[0:0];
  _RAND_400 = {1{`RANDOM}};
  dataArray_8_5_cachedata_MPORT_en_pipe_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dataArray_8_5_cachedata_MPORT_addr_pipe_0 = _RAND_401[0:0];
  _RAND_403 = {1{`RANDOM}};
  dataArray_8_6_cachedata_MPORT_en_pipe_0 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dataArray_8_6_cachedata_MPORT_addr_pipe_0 = _RAND_404[0:0];
  _RAND_406 = {1{`RANDOM}};
  dataArray_8_7_cachedata_MPORT_en_pipe_0 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dataArray_8_7_cachedata_MPORT_addr_pipe_0 = _RAND_407[0:0];
  _RAND_409 = {1{`RANDOM}};
  dataArray_8_8_cachedata_MPORT_en_pipe_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dataArray_8_8_cachedata_MPORT_addr_pipe_0 = _RAND_410[0:0];
  _RAND_412 = {1{`RANDOM}};
  dataArray_8_9_cachedata_MPORT_en_pipe_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dataArray_8_9_cachedata_MPORT_addr_pipe_0 = _RAND_413[0:0];
  _RAND_415 = {1{`RANDOM}};
  dataArray_8_10_cachedata_MPORT_en_pipe_0 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dataArray_8_10_cachedata_MPORT_addr_pipe_0 = _RAND_416[0:0];
  _RAND_418 = {1{`RANDOM}};
  dataArray_8_11_cachedata_MPORT_en_pipe_0 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dataArray_8_11_cachedata_MPORT_addr_pipe_0 = _RAND_419[0:0];
  _RAND_421 = {1{`RANDOM}};
  dataArray_8_12_cachedata_MPORT_en_pipe_0 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dataArray_8_12_cachedata_MPORT_addr_pipe_0 = _RAND_422[0:0];
  _RAND_424 = {1{`RANDOM}};
  dataArray_8_13_cachedata_MPORT_en_pipe_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dataArray_8_13_cachedata_MPORT_addr_pipe_0 = _RAND_425[0:0];
  _RAND_427 = {1{`RANDOM}};
  dataArray_8_14_cachedata_MPORT_en_pipe_0 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dataArray_8_14_cachedata_MPORT_addr_pipe_0 = _RAND_428[0:0];
  _RAND_430 = {1{`RANDOM}};
  dataArray_8_15_cachedata_MPORT_en_pipe_0 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dataArray_8_15_cachedata_MPORT_addr_pipe_0 = _RAND_431[0:0];
  _RAND_433 = {1{`RANDOM}};
  dataArray_9_0_cachedata_MPORT_en_pipe_0 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dataArray_9_0_cachedata_MPORT_addr_pipe_0 = _RAND_434[0:0];
  _RAND_436 = {1{`RANDOM}};
  dataArray_9_1_cachedata_MPORT_en_pipe_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dataArray_9_1_cachedata_MPORT_addr_pipe_0 = _RAND_437[0:0];
  _RAND_439 = {1{`RANDOM}};
  dataArray_9_2_cachedata_MPORT_en_pipe_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dataArray_9_2_cachedata_MPORT_addr_pipe_0 = _RAND_440[0:0];
  _RAND_442 = {1{`RANDOM}};
  dataArray_9_3_cachedata_MPORT_en_pipe_0 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dataArray_9_3_cachedata_MPORT_addr_pipe_0 = _RAND_443[0:0];
  _RAND_445 = {1{`RANDOM}};
  dataArray_9_4_cachedata_MPORT_en_pipe_0 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dataArray_9_4_cachedata_MPORT_addr_pipe_0 = _RAND_446[0:0];
  _RAND_448 = {1{`RANDOM}};
  dataArray_9_5_cachedata_MPORT_en_pipe_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dataArray_9_5_cachedata_MPORT_addr_pipe_0 = _RAND_449[0:0];
  _RAND_451 = {1{`RANDOM}};
  dataArray_9_6_cachedata_MPORT_en_pipe_0 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dataArray_9_6_cachedata_MPORT_addr_pipe_0 = _RAND_452[0:0];
  _RAND_454 = {1{`RANDOM}};
  dataArray_9_7_cachedata_MPORT_en_pipe_0 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dataArray_9_7_cachedata_MPORT_addr_pipe_0 = _RAND_455[0:0];
  _RAND_457 = {1{`RANDOM}};
  dataArray_9_8_cachedata_MPORT_en_pipe_0 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dataArray_9_8_cachedata_MPORT_addr_pipe_0 = _RAND_458[0:0];
  _RAND_460 = {1{`RANDOM}};
  dataArray_9_9_cachedata_MPORT_en_pipe_0 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dataArray_9_9_cachedata_MPORT_addr_pipe_0 = _RAND_461[0:0];
  _RAND_463 = {1{`RANDOM}};
  dataArray_9_10_cachedata_MPORT_en_pipe_0 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dataArray_9_10_cachedata_MPORT_addr_pipe_0 = _RAND_464[0:0];
  _RAND_466 = {1{`RANDOM}};
  dataArray_9_11_cachedata_MPORT_en_pipe_0 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dataArray_9_11_cachedata_MPORT_addr_pipe_0 = _RAND_467[0:0];
  _RAND_469 = {1{`RANDOM}};
  dataArray_9_12_cachedata_MPORT_en_pipe_0 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dataArray_9_12_cachedata_MPORT_addr_pipe_0 = _RAND_470[0:0];
  _RAND_472 = {1{`RANDOM}};
  dataArray_9_13_cachedata_MPORT_en_pipe_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dataArray_9_13_cachedata_MPORT_addr_pipe_0 = _RAND_473[0:0];
  _RAND_475 = {1{`RANDOM}};
  dataArray_9_14_cachedata_MPORT_en_pipe_0 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dataArray_9_14_cachedata_MPORT_addr_pipe_0 = _RAND_476[0:0];
  _RAND_478 = {1{`RANDOM}};
  dataArray_9_15_cachedata_MPORT_en_pipe_0 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dataArray_9_15_cachedata_MPORT_addr_pipe_0 = _RAND_479[0:0];
  _RAND_481 = {1{`RANDOM}};
  dataArray_10_0_cachedata_MPORT_en_pipe_0 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dataArray_10_0_cachedata_MPORT_addr_pipe_0 = _RAND_482[0:0];
  _RAND_484 = {1{`RANDOM}};
  dataArray_10_1_cachedata_MPORT_en_pipe_0 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dataArray_10_1_cachedata_MPORT_addr_pipe_0 = _RAND_485[0:0];
  _RAND_487 = {1{`RANDOM}};
  dataArray_10_2_cachedata_MPORT_en_pipe_0 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dataArray_10_2_cachedata_MPORT_addr_pipe_0 = _RAND_488[0:0];
  _RAND_490 = {1{`RANDOM}};
  dataArray_10_3_cachedata_MPORT_en_pipe_0 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dataArray_10_3_cachedata_MPORT_addr_pipe_0 = _RAND_491[0:0];
  _RAND_493 = {1{`RANDOM}};
  dataArray_10_4_cachedata_MPORT_en_pipe_0 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dataArray_10_4_cachedata_MPORT_addr_pipe_0 = _RAND_494[0:0];
  _RAND_496 = {1{`RANDOM}};
  dataArray_10_5_cachedata_MPORT_en_pipe_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dataArray_10_5_cachedata_MPORT_addr_pipe_0 = _RAND_497[0:0];
  _RAND_499 = {1{`RANDOM}};
  dataArray_10_6_cachedata_MPORT_en_pipe_0 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dataArray_10_6_cachedata_MPORT_addr_pipe_0 = _RAND_500[0:0];
  _RAND_502 = {1{`RANDOM}};
  dataArray_10_7_cachedata_MPORT_en_pipe_0 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dataArray_10_7_cachedata_MPORT_addr_pipe_0 = _RAND_503[0:0];
  _RAND_505 = {1{`RANDOM}};
  dataArray_10_8_cachedata_MPORT_en_pipe_0 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dataArray_10_8_cachedata_MPORT_addr_pipe_0 = _RAND_506[0:0];
  _RAND_508 = {1{`RANDOM}};
  dataArray_10_9_cachedata_MPORT_en_pipe_0 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dataArray_10_9_cachedata_MPORT_addr_pipe_0 = _RAND_509[0:0];
  _RAND_511 = {1{`RANDOM}};
  dataArray_10_10_cachedata_MPORT_en_pipe_0 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dataArray_10_10_cachedata_MPORT_addr_pipe_0 = _RAND_512[0:0];
  _RAND_514 = {1{`RANDOM}};
  dataArray_10_11_cachedata_MPORT_en_pipe_0 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dataArray_10_11_cachedata_MPORT_addr_pipe_0 = _RAND_515[0:0];
  _RAND_517 = {1{`RANDOM}};
  dataArray_10_12_cachedata_MPORT_en_pipe_0 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  dataArray_10_12_cachedata_MPORT_addr_pipe_0 = _RAND_518[0:0];
  _RAND_520 = {1{`RANDOM}};
  dataArray_10_13_cachedata_MPORT_en_pipe_0 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  dataArray_10_13_cachedata_MPORT_addr_pipe_0 = _RAND_521[0:0];
  _RAND_523 = {1{`RANDOM}};
  dataArray_10_14_cachedata_MPORT_en_pipe_0 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  dataArray_10_14_cachedata_MPORT_addr_pipe_0 = _RAND_524[0:0];
  _RAND_526 = {1{`RANDOM}};
  dataArray_10_15_cachedata_MPORT_en_pipe_0 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  dataArray_10_15_cachedata_MPORT_addr_pipe_0 = _RAND_527[0:0];
  _RAND_529 = {1{`RANDOM}};
  dataArray_11_0_cachedata_MPORT_en_pipe_0 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dataArray_11_0_cachedata_MPORT_addr_pipe_0 = _RAND_530[0:0];
  _RAND_532 = {1{`RANDOM}};
  dataArray_11_1_cachedata_MPORT_en_pipe_0 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dataArray_11_1_cachedata_MPORT_addr_pipe_0 = _RAND_533[0:0];
  _RAND_535 = {1{`RANDOM}};
  dataArray_11_2_cachedata_MPORT_en_pipe_0 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  dataArray_11_2_cachedata_MPORT_addr_pipe_0 = _RAND_536[0:0];
  _RAND_538 = {1{`RANDOM}};
  dataArray_11_3_cachedata_MPORT_en_pipe_0 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  dataArray_11_3_cachedata_MPORT_addr_pipe_0 = _RAND_539[0:0];
  _RAND_541 = {1{`RANDOM}};
  dataArray_11_4_cachedata_MPORT_en_pipe_0 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  dataArray_11_4_cachedata_MPORT_addr_pipe_0 = _RAND_542[0:0];
  _RAND_544 = {1{`RANDOM}};
  dataArray_11_5_cachedata_MPORT_en_pipe_0 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  dataArray_11_5_cachedata_MPORT_addr_pipe_0 = _RAND_545[0:0];
  _RAND_547 = {1{`RANDOM}};
  dataArray_11_6_cachedata_MPORT_en_pipe_0 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  dataArray_11_6_cachedata_MPORT_addr_pipe_0 = _RAND_548[0:0];
  _RAND_550 = {1{`RANDOM}};
  dataArray_11_7_cachedata_MPORT_en_pipe_0 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  dataArray_11_7_cachedata_MPORT_addr_pipe_0 = _RAND_551[0:0];
  _RAND_553 = {1{`RANDOM}};
  dataArray_11_8_cachedata_MPORT_en_pipe_0 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dataArray_11_8_cachedata_MPORT_addr_pipe_0 = _RAND_554[0:0];
  _RAND_556 = {1{`RANDOM}};
  dataArray_11_9_cachedata_MPORT_en_pipe_0 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  dataArray_11_9_cachedata_MPORT_addr_pipe_0 = _RAND_557[0:0];
  _RAND_559 = {1{`RANDOM}};
  dataArray_11_10_cachedata_MPORT_en_pipe_0 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  dataArray_11_10_cachedata_MPORT_addr_pipe_0 = _RAND_560[0:0];
  _RAND_562 = {1{`RANDOM}};
  dataArray_11_11_cachedata_MPORT_en_pipe_0 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  dataArray_11_11_cachedata_MPORT_addr_pipe_0 = _RAND_563[0:0];
  _RAND_565 = {1{`RANDOM}};
  dataArray_11_12_cachedata_MPORT_en_pipe_0 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  dataArray_11_12_cachedata_MPORT_addr_pipe_0 = _RAND_566[0:0];
  _RAND_568 = {1{`RANDOM}};
  dataArray_11_13_cachedata_MPORT_en_pipe_0 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  dataArray_11_13_cachedata_MPORT_addr_pipe_0 = _RAND_569[0:0];
  _RAND_571 = {1{`RANDOM}};
  dataArray_11_14_cachedata_MPORT_en_pipe_0 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  dataArray_11_14_cachedata_MPORT_addr_pipe_0 = _RAND_572[0:0];
  _RAND_574 = {1{`RANDOM}};
  dataArray_11_15_cachedata_MPORT_en_pipe_0 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  dataArray_11_15_cachedata_MPORT_addr_pipe_0 = _RAND_575[0:0];
  _RAND_577 = {1{`RANDOM}};
  dataArray_12_0_cachedata_MPORT_en_pipe_0 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  dataArray_12_0_cachedata_MPORT_addr_pipe_0 = _RAND_578[0:0];
  _RAND_580 = {1{`RANDOM}};
  dataArray_12_1_cachedata_MPORT_en_pipe_0 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  dataArray_12_1_cachedata_MPORT_addr_pipe_0 = _RAND_581[0:0];
  _RAND_583 = {1{`RANDOM}};
  dataArray_12_2_cachedata_MPORT_en_pipe_0 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  dataArray_12_2_cachedata_MPORT_addr_pipe_0 = _RAND_584[0:0];
  _RAND_586 = {1{`RANDOM}};
  dataArray_12_3_cachedata_MPORT_en_pipe_0 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  dataArray_12_3_cachedata_MPORT_addr_pipe_0 = _RAND_587[0:0];
  _RAND_589 = {1{`RANDOM}};
  dataArray_12_4_cachedata_MPORT_en_pipe_0 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  dataArray_12_4_cachedata_MPORT_addr_pipe_0 = _RAND_590[0:0];
  _RAND_592 = {1{`RANDOM}};
  dataArray_12_5_cachedata_MPORT_en_pipe_0 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  dataArray_12_5_cachedata_MPORT_addr_pipe_0 = _RAND_593[0:0];
  _RAND_595 = {1{`RANDOM}};
  dataArray_12_6_cachedata_MPORT_en_pipe_0 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  dataArray_12_6_cachedata_MPORT_addr_pipe_0 = _RAND_596[0:0];
  _RAND_598 = {1{`RANDOM}};
  dataArray_12_7_cachedata_MPORT_en_pipe_0 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  dataArray_12_7_cachedata_MPORT_addr_pipe_0 = _RAND_599[0:0];
  _RAND_601 = {1{`RANDOM}};
  dataArray_12_8_cachedata_MPORT_en_pipe_0 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  dataArray_12_8_cachedata_MPORT_addr_pipe_0 = _RAND_602[0:0];
  _RAND_604 = {1{`RANDOM}};
  dataArray_12_9_cachedata_MPORT_en_pipe_0 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  dataArray_12_9_cachedata_MPORT_addr_pipe_0 = _RAND_605[0:0];
  _RAND_607 = {1{`RANDOM}};
  dataArray_12_10_cachedata_MPORT_en_pipe_0 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  dataArray_12_10_cachedata_MPORT_addr_pipe_0 = _RAND_608[0:0];
  _RAND_610 = {1{`RANDOM}};
  dataArray_12_11_cachedata_MPORT_en_pipe_0 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  dataArray_12_11_cachedata_MPORT_addr_pipe_0 = _RAND_611[0:0];
  _RAND_613 = {1{`RANDOM}};
  dataArray_12_12_cachedata_MPORT_en_pipe_0 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  dataArray_12_12_cachedata_MPORT_addr_pipe_0 = _RAND_614[0:0];
  _RAND_616 = {1{`RANDOM}};
  dataArray_12_13_cachedata_MPORT_en_pipe_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  dataArray_12_13_cachedata_MPORT_addr_pipe_0 = _RAND_617[0:0];
  _RAND_619 = {1{`RANDOM}};
  dataArray_12_14_cachedata_MPORT_en_pipe_0 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  dataArray_12_14_cachedata_MPORT_addr_pipe_0 = _RAND_620[0:0];
  _RAND_622 = {1{`RANDOM}};
  dataArray_12_15_cachedata_MPORT_en_pipe_0 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  dataArray_12_15_cachedata_MPORT_addr_pipe_0 = _RAND_623[0:0];
  _RAND_625 = {1{`RANDOM}};
  dataArray_13_0_cachedata_MPORT_en_pipe_0 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  dataArray_13_0_cachedata_MPORT_addr_pipe_0 = _RAND_626[0:0];
  _RAND_628 = {1{`RANDOM}};
  dataArray_13_1_cachedata_MPORT_en_pipe_0 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  dataArray_13_1_cachedata_MPORT_addr_pipe_0 = _RAND_629[0:0];
  _RAND_631 = {1{`RANDOM}};
  dataArray_13_2_cachedata_MPORT_en_pipe_0 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  dataArray_13_2_cachedata_MPORT_addr_pipe_0 = _RAND_632[0:0];
  _RAND_634 = {1{`RANDOM}};
  dataArray_13_3_cachedata_MPORT_en_pipe_0 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  dataArray_13_3_cachedata_MPORT_addr_pipe_0 = _RAND_635[0:0];
  _RAND_637 = {1{`RANDOM}};
  dataArray_13_4_cachedata_MPORT_en_pipe_0 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  dataArray_13_4_cachedata_MPORT_addr_pipe_0 = _RAND_638[0:0];
  _RAND_640 = {1{`RANDOM}};
  dataArray_13_5_cachedata_MPORT_en_pipe_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  dataArray_13_5_cachedata_MPORT_addr_pipe_0 = _RAND_641[0:0];
  _RAND_643 = {1{`RANDOM}};
  dataArray_13_6_cachedata_MPORT_en_pipe_0 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  dataArray_13_6_cachedata_MPORT_addr_pipe_0 = _RAND_644[0:0];
  _RAND_646 = {1{`RANDOM}};
  dataArray_13_7_cachedata_MPORT_en_pipe_0 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  dataArray_13_7_cachedata_MPORT_addr_pipe_0 = _RAND_647[0:0];
  _RAND_649 = {1{`RANDOM}};
  dataArray_13_8_cachedata_MPORT_en_pipe_0 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  dataArray_13_8_cachedata_MPORT_addr_pipe_0 = _RAND_650[0:0];
  _RAND_652 = {1{`RANDOM}};
  dataArray_13_9_cachedata_MPORT_en_pipe_0 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  dataArray_13_9_cachedata_MPORT_addr_pipe_0 = _RAND_653[0:0];
  _RAND_655 = {1{`RANDOM}};
  dataArray_13_10_cachedata_MPORT_en_pipe_0 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  dataArray_13_10_cachedata_MPORT_addr_pipe_0 = _RAND_656[0:0];
  _RAND_658 = {1{`RANDOM}};
  dataArray_13_11_cachedata_MPORT_en_pipe_0 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  dataArray_13_11_cachedata_MPORT_addr_pipe_0 = _RAND_659[0:0];
  _RAND_661 = {1{`RANDOM}};
  dataArray_13_12_cachedata_MPORT_en_pipe_0 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  dataArray_13_12_cachedata_MPORT_addr_pipe_0 = _RAND_662[0:0];
  _RAND_664 = {1{`RANDOM}};
  dataArray_13_13_cachedata_MPORT_en_pipe_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  dataArray_13_13_cachedata_MPORT_addr_pipe_0 = _RAND_665[0:0];
  _RAND_667 = {1{`RANDOM}};
  dataArray_13_14_cachedata_MPORT_en_pipe_0 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  dataArray_13_14_cachedata_MPORT_addr_pipe_0 = _RAND_668[0:0];
  _RAND_670 = {1{`RANDOM}};
  dataArray_13_15_cachedata_MPORT_en_pipe_0 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  dataArray_13_15_cachedata_MPORT_addr_pipe_0 = _RAND_671[0:0];
  _RAND_673 = {1{`RANDOM}};
  dataArray_14_0_cachedata_MPORT_en_pipe_0 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  dataArray_14_0_cachedata_MPORT_addr_pipe_0 = _RAND_674[0:0];
  _RAND_676 = {1{`RANDOM}};
  dataArray_14_1_cachedata_MPORT_en_pipe_0 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  dataArray_14_1_cachedata_MPORT_addr_pipe_0 = _RAND_677[0:0];
  _RAND_679 = {1{`RANDOM}};
  dataArray_14_2_cachedata_MPORT_en_pipe_0 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  dataArray_14_2_cachedata_MPORT_addr_pipe_0 = _RAND_680[0:0];
  _RAND_682 = {1{`RANDOM}};
  dataArray_14_3_cachedata_MPORT_en_pipe_0 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  dataArray_14_3_cachedata_MPORT_addr_pipe_0 = _RAND_683[0:0];
  _RAND_685 = {1{`RANDOM}};
  dataArray_14_4_cachedata_MPORT_en_pipe_0 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  dataArray_14_4_cachedata_MPORT_addr_pipe_0 = _RAND_686[0:0];
  _RAND_688 = {1{`RANDOM}};
  dataArray_14_5_cachedata_MPORT_en_pipe_0 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  dataArray_14_5_cachedata_MPORT_addr_pipe_0 = _RAND_689[0:0];
  _RAND_691 = {1{`RANDOM}};
  dataArray_14_6_cachedata_MPORT_en_pipe_0 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  dataArray_14_6_cachedata_MPORT_addr_pipe_0 = _RAND_692[0:0];
  _RAND_694 = {1{`RANDOM}};
  dataArray_14_7_cachedata_MPORT_en_pipe_0 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  dataArray_14_7_cachedata_MPORT_addr_pipe_0 = _RAND_695[0:0];
  _RAND_697 = {1{`RANDOM}};
  dataArray_14_8_cachedata_MPORT_en_pipe_0 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  dataArray_14_8_cachedata_MPORT_addr_pipe_0 = _RAND_698[0:0];
  _RAND_700 = {1{`RANDOM}};
  dataArray_14_9_cachedata_MPORT_en_pipe_0 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  dataArray_14_9_cachedata_MPORT_addr_pipe_0 = _RAND_701[0:0];
  _RAND_703 = {1{`RANDOM}};
  dataArray_14_10_cachedata_MPORT_en_pipe_0 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  dataArray_14_10_cachedata_MPORT_addr_pipe_0 = _RAND_704[0:0];
  _RAND_706 = {1{`RANDOM}};
  dataArray_14_11_cachedata_MPORT_en_pipe_0 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  dataArray_14_11_cachedata_MPORT_addr_pipe_0 = _RAND_707[0:0];
  _RAND_709 = {1{`RANDOM}};
  dataArray_14_12_cachedata_MPORT_en_pipe_0 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  dataArray_14_12_cachedata_MPORT_addr_pipe_0 = _RAND_710[0:0];
  _RAND_712 = {1{`RANDOM}};
  dataArray_14_13_cachedata_MPORT_en_pipe_0 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  dataArray_14_13_cachedata_MPORT_addr_pipe_0 = _RAND_713[0:0];
  _RAND_715 = {1{`RANDOM}};
  dataArray_14_14_cachedata_MPORT_en_pipe_0 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  dataArray_14_14_cachedata_MPORT_addr_pipe_0 = _RAND_716[0:0];
  _RAND_718 = {1{`RANDOM}};
  dataArray_14_15_cachedata_MPORT_en_pipe_0 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  dataArray_14_15_cachedata_MPORT_addr_pipe_0 = _RAND_719[0:0];
  _RAND_721 = {1{`RANDOM}};
  dataArray_15_0_cachedata_MPORT_en_pipe_0 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  dataArray_15_0_cachedata_MPORT_addr_pipe_0 = _RAND_722[0:0];
  _RAND_724 = {1{`RANDOM}};
  dataArray_15_1_cachedata_MPORT_en_pipe_0 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  dataArray_15_1_cachedata_MPORT_addr_pipe_0 = _RAND_725[0:0];
  _RAND_727 = {1{`RANDOM}};
  dataArray_15_2_cachedata_MPORT_en_pipe_0 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  dataArray_15_2_cachedata_MPORT_addr_pipe_0 = _RAND_728[0:0];
  _RAND_730 = {1{`RANDOM}};
  dataArray_15_3_cachedata_MPORT_en_pipe_0 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  dataArray_15_3_cachedata_MPORT_addr_pipe_0 = _RAND_731[0:0];
  _RAND_733 = {1{`RANDOM}};
  dataArray_15_4_cachedata_MPORT_en_pipe_0 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  dataArray_15_4_cachedata_MPORT_addr_pipe_0 = _RAND_734[0:0];
  _RAND_736 = {1{`RANDOM}};
  dataArray_15_5_cachedata_MPORT_en_pipe_0 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  dataArray_15_5_cachedata_MPORT_addr_pipe_0 = _RAND_737[0:0];
  _RAND_739 = {1{`RANDOM}};
  dataArray_15_6_cachedata_MPORT_en_pipe_0 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  dataArray_15_6_cachedata_MPORT_addr_pipe_0 = _RAND_740[0:0];
  _RAND_742 = {1{`RANDOM}};
  dataArray_15_7_cachedata_MPORT_en_pipe_0 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  dataArray_15_7_cachedata_MPORT_addr_pipe_0 = _RAND_743[0:0];
  _RAND_745 = {1{`RANDOM}};
  dataArray_15_8_cachedata_MPORT_en_pipe_0 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  dataArray_15_8_cachedata_MPORT_addr_pipe_0 = _RAND_746[0:0];
  _RAND_748 = {1{`RANDOM}};
  dataArray_15_9_cachedata_MPORT_en_pipe_0 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  dataArray_15_9_cachedata_MPORT_addr_pipe_0 = _RAND_749[0:0];
  _RAND_751 = {1{`RANDOM}};
  dataArray_15_10_cachedata_MPORT_en_pipe_0 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  dataArray_15_10_cachedata_MPORT_addr_pipe_0 = _RAND_752[0:0];
  _RAND_754 = {1{`RANDOM}};
  dataArray_15_11_cachedata_MPORT_en_pipe_0 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  dataArray_15_11_cachedata_MPORT_addr_pipe_0 = _RAND_755[0:0];
  _RAND_757 = {1{`RANDOM}};
  dataArray_15_12_cachedata_MPORT_en_pipe_0 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  dataArray_15_12_cachedata_MPORT_addr_pipe_0 = _RAND_758[0:0];
  _RAND_760 = {1{`RANDOM}};
  dataArray_15_13_cachedata_MPORT_en_pipe_0 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  dataArray_15_13_cachedata_MPORT_addr_pipe_0 = _RAND_761[0:0];
  _RAND_763 = {1{`RANDOM}};
  dataArray_15_14_cachedata_MPORT_en_pipe_0 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  dataArray_15_14_cachedata_MPORT_addr_pipe_0 = _RAND_764[0:0];
  _RAND_766 = {1{`RANDOM}};
  dataArray_15_15_cachedata_MPORT_en_pipe_0 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  dataArray_15_15_cachedata_MPORT_addr_pipe_0 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  replace_set = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  random_num = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  tagArray_0_0 = _RAND_770[21:0];
  _RAND_771 = {1{`RANDOM}};
  tagArray_0_1 = _RAND_771[21:0];
  _RAND_772 = {1{`RANDOM}};
  tagArray_0_2 = _RAND_772[21:0];
  _RAND_773 = {1{`RANDOM}};
  tagArray_0_3 = _RAND_773[21:0];
  _RAND_774 = {1{`RANDOM}};
  tagArray_0_4 = _RAND_774[21:0];
  _RAND_775 = {1{`RANDOM}};
  tagArray_0_5 = _RAND_775[21:0];
  _RAND_776 = {1{`RANDOM}};
  tagArray_0_6 = _RAND_776[21:0];
  _RAND_777 = {1{`RANDOM}};
  tagArray_0_7 = _RAND_777[21:0];
  _RAND_778 = {1{`RANDOM}};
  tagArray_0_8 = _RAND_778[21:0];
  _RAND_779 = {1{`RANDOM}};
  tagArray_0_9 = _RAND_779[21:0];
  _RAND_780 = {1{`RANDOM}};
  tagArray_0_10 = _RAND_780[21:0];
  _RAND_781 = {1{`RANDOM}};
  tagArray_0_11 = _RAND_781[21:0];
  _RAND_782 = {1{`RANDOM}};
  tagArray_0_12 = _RAND_782[21:0];
  _RAND_783 = {1{`RANDOM}};
  tagArray_0_13 = _RAND_783[21:0];
  _RAND_784 = {1{`RANDOM}};
  tagArray_0_14 = _RAND_784[21:0];
  _RAND_785 = {1{`RANDOM}};
  tagArray_0_15 = _RAND_785[21:0];
  _RAND_786 = {1{`RANDOM}};
  tagArray_1_0 = _RAND_786[21:0];
  _RAND_787 = {1{`RANDOM}};
  tagArray_1_1 = _RAND_787[21:0];
  _RAND_788 = {1{`RANDOM}};
  tagArray_1_2 = _RAND_788[21:0];
  _RAND_789 = {1{`RANDOM}};
  tagArray_1_3 = _RAND_789[21:0];
  _RAND_790 = {1{`RANDOM}};
  tagArray_1_4 = _RAND_790[21:0];
  _RAND_791 = {1{`RANDOM}};
  tagArray_1_5 = _RAND_791[21:0];
  _RAND_792 = {1{`RANDOM}};
  tagArray_1_6 = _RAND_792[21:0];
  _RAND_793 = {1{`RANDOM}};
  tagArray_1_7 = _RAND_793[21:0];
  _RAND_794 = {1{`RANDOM}};
  tagArray_1_8 = _RAND_794[21:0];
  _RAND_795 = {1{`RANDOM}};
  tagArray_1_9 = _RAND_795[21:0];
  _RAND_796 = {1{`RANDOM}};
  tagArray_1_10 = _RAND_796[21:0];
  _RAND_797 = {1{`RANDOM}};
  tagArray_1_11 = _RAND_797[21:0];
  _RAND_798 = {1{`RANDOM}};
  tagArray_1_12 = _RAND_798[21:0];
  _RAND_799 = {1{`RANDOM}};
  tagArray_1_13 = _RAND_799[21:0];
  _RAND_800 = {1{`RANDOM}};
  tagArray_1_14 = _RAND_800[21:0];
  _RAND_801 = {1{`RANDOM}};
  tagArray_1_15 = _RAND_801[21:0];
  _RAND_802 = {1{`RANDOM}};
  validArray_0_0 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  validArray_0_1 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  validArray_0_2 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  validArray_0_3 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  validArray_0_4 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  validArray_0_5 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  validArray_0_6 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  validArray_0_7 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  validArray_0_8 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  validArray_0_9 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  validArray_0_10 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  validArray_0_11 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  validArray_0_12 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  validArray_0_13 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  validArray_0_14 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  validArray_0_15 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  validArray_1_0 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  validArray_1_1 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  validArray_1_2 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  validArray_1_3 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  validArray_1_4 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  validArray_1_5 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  validArray_1_6 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  validArray_1_7 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  validArray_1_8 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  validArray_1_9 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  validArray_1_10 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  validArray_1_11 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  validArray_1_12 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  validArray_1_13 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  validArray_1_14 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  validArray_1_15 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  off = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  state_cache = _RAND_835[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAM_axi(
  input         clock,
  input         reset,
  output        axi_ar_ready,
  input         axi_ar_valid,
  input  [31:0] axi_ar_bits_addr,
  input  [7:0]  axi_ar_bits_len,
  input         axi_r_ready,
  output        axi_r_valid,
  output [31:0] axi_r_bits_data,
  output        axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  RamBB_i1_clock; // @[sram_Axi.scala 65:26]
  wire [31:0] RamBB_i1_addr; // @[sram_Axi.scala 65:26]
  wire  RamBB_i1_mem_wen; // @[sram_Axi.scala 65:26]
  wire  RamBB_i1_valid; // @[sram_Axi.scala 65:26]
  wire [31:0] RamBB_i1_wdata; // @[sram_Axi.scala 65:26]
  wire [3:0] RamBB_i1_wmask; // @[sram_Axi.scala 65:26]
  wire [31:0] RamBB_i1_rdata; // @[sram_Axi.scala 65:26]
  reg  delay; // @[sram_Axi.scala 22:24]
  reg [7:0] reg_AxLen; // @[sram_Axi.scala 25:28]
  reg [31:0] reg_addr; // @[sram_Axi.scala 26:28]
  reg [1:0] reg_burst; // @[sram_Axi.scala 27:28]
  reg [1:0] state_sram; // @[sram_Axi.scala 31:29]
  wire  _T_1 = axi_ar_ready & axi_ar_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_sram_T_1 = reg_AxLen == 8'h0 ? 2'h3 : 2'h2; // @[sram_Axi.scala 47:34]
  wire  _T_4 = 2'h2 == state_sram; // @[sram_Axi.scala 32:25]
  wire [1:0] _state_sram_T_3 = reg_AxLen == 8'h1 ? 2'h3 : 2'h2; // @[sram_Axi.scala 54:31]
  wire  _reg_AxLen_T = axi_r_ready & axi_r_valid; // @[Decoupled.scala 51:35]
  wire [7:0] _reg_AxLen_T_2 = reg_AxLen - 8'h1; // @[sram_Axi.scala 55:53]
  wire [7:0] _reg_AxLen_T_3 = _reg_AxLen_T ? _reg_AxLen_T_2 : reg_AxLen; // @[sram_Axi.scala 55:31]
  wire [31:0] _reg_addr_T_2 = reg_addr + 32'h4; // @[sram_Axi.scala 57:53]
  wire [31:0] _reg_addr_T_3 = _reg_AxLen_T ? _reg_addr_T_2 : reg_addr; // @[sram_Axi.scala 57:30]
  wire [31:0] _reg_addr_T_5 = 2'h1 == reg_burst ? _reg_addr_T_3 : reg_addr; // @[Mux.scala 81:58]
  wire  _T_5 = 2'h3 == state_sram; // @[sram_Axi.scala 32:25]
  wire [1:0] _GEN_5 = 2'h3 == state_sram ? 2'h0 : state_sram; // @[sram_Axi.scala 32:25 61:24 31:29]
  RamBB RamBB_i1 ( // @[sram_Axi.scala 65:26]
    .clock(RamBB_i1_clock),
    .addr(RamBB_i1_addr),
    .mem_wen(RamBB_i1_mem_wen),
    .valid(RamBB_i1_valid),
    .wdata(RamBB_i1_wdata),
    .wmask(RamBB_i1_wmask),
    .rdata(RamBB_i1_rdata)
  );
  assign axi_ar_ready = 2'h0 == state_sram; // @[Mux.scala 81:61]
  assign axi_r_valid = _T_5 | _T_4; // @[Mux.scala 81:58]
  assign axi_r_bits_data = RamBB_i1_rdata; // @[sram_Axi.scala 78:21]
  assign axi_r_bits_last = state_sram == 2'h3; // @[sram_Axi.scala 80:39]
  assign RamBB_i1_clock = clock; // @[sram_Axi.scala 66:25]
  assign RamBB_i1_addr = reg_addr; // @[sram_Axi.scala 67:25]
  assign RamBB_i1_mem_wen = 1'h0; // @[sram_Axi.scala 68:25]
  assign RamBB_i1_valid = _T_5 | _T_4; // @[Mux.scala 81:58]
  assign RamBB_i1_wdata = 32'h0; // @[sram_Axi.scala 72:25]
  assign RamBB_i1_wmask = 4'h0; // @[sram_Axi.scala 73:25]
  always @(posedge clock) begin
    if (reset) begin // @[sram_Axi.scala 22:24]
      delay <= 1'h0; // @[sram_Axi.scala 22:24]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      delay <= 1'h0; // @[sram_Axi.scala 34:19]
    end else if (2'h1 == state_sram) begin // @[sram_Axi.scala 32:25]
      delay <= delay - 1'h1; // @[sram_Axi.scala 51:19]
    end
    if (reset) begin // @[sram_Axi.scala 25:28]
      reg_AxLen <= 8'h0; // @[sram_Axi.scala 25:28]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        reg_AxLen <= axi_ar_bits_len; // @[sram_Axi.scala 38:28]
      end
    end else if (!(2'h1 == state_sram)) begin // @[sram_Axi.scala 32:25]
      if (2'h2 == state_sram) begin // @[sram_Axi.scala 32:25]
        reg_AxLen <= _reg_AxLen_T_3; // @[sram_Axi.scala 55:25]
      end
    end
    if (reset) begin // @[sram_Axi.scala 26:28]
      reg_addr <= 32'h0; // @[sram_Axi.scala 26:28]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        reg_addr <= axi_ar_bits_addr; // @[sram_Axi.scala 39:28]
      end
    end else if (!(2'h1 == state_sram)) begin // @[sram_Axi.scala 32:25]
      if (2'h2 == state_sram) begin // @[sram_Axi.scala 32:25]
        reg_addr <= _reg_addr_T_5; // @[sram_Axi.scala 56:25]
      end
    end
    if (reset) begin // @[sram_Axi.scala 27:28]
      reg_burst <= 2'h3; // @[sram_Axi.scala 27:28]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        reg_burst <= 2'h1; // @[sram_Axi.scala 40:28]
      end
    end
    if (reset) begin // @[sram_Axi.scala 31:29]
      state_sram <= 2'h0; // @[sram_Axi.scala 31:29]
    end else if (2'h0 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (_T_1) begin // @[sram_Axi.scala 36:32]
        state_sram <= 2'h1; // @[sram_Axi.scala 37:28]
      end else begin
        state_sram <= 2'h0; // @[sram_Axi.scala 42:28]
      end
    end else if (2'h1 == state_sram) begin // @[sram_Axi.scala 32:25]
      if (~delay) begin // @[sram_Axi.scala 46:34]
        state_sram <= _state_sram_T_1; // @[sram_Axi.scala 47:28]
      end else begin
        state_sram <= 2'h1; // @[sram_Axi.scala 49:28]
      end
    end else if (2'h2 == state_sram) begin // @[sram_Axi.scala 32:25]
      state_sram <= _state_sram_T_3; // @[sram_Axi.scala 54:25]
    end else begin
      state_sram <= _GEN_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_AxLen = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  reg_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_burst = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  state_sram = _RAND_4[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAM(
  input         clock,
  input         reset,
  output        axi_ar_ready,
  input         axi_ar_valid,
  input  [31:0] axi_ar_bits_addr,
  input         axi_r_ready,
  output        axi_r_valid,
  output [31:0] axi_r_bits_data,
  output        axi_aw_ready,
  input         axi_aw_valid,
  input  [31:0] axi_aw_bits_addr,
  output        axi_w_ready,
  input         axi_w_valid,
  input  [31:0] axi_w_bits_data,
  input  [3:0]  axi_w_bits_strb,
  input         axi_b_ready,
  output        axi_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RamBB_i1_clock; // @[sram_AxiLite.scala 77:26]
  wire [31:0] RamBB_i1_addr; // @[sram_AxiLite.scala 77:26]
  wire  RamBB_i1_mem_wen; // @[sram_AxiLite.scala 77:26]
  wire  RamBB_i1_valid; // @[sram_AxiLite.scala 77:26]
  wire [31:0] RamBB_i1_wdata; // @[sram_AxiLite.scala 77:26]
  wire [3:0] RamBB_i1_wmask; // @[sram_AxiLite.scala 77:26]
  wire [31:0] RamBB_i1_rdata; // @[sram_AxiLite.scala 77:26]
  reg  delay; // @[sram_AxiLite.scala 42:24]
  reg [2:0] state; // @[sram_AxiLite.scala 46:24]
  wire  _T_1 = axi_ar_ready & axi_ar_valid; // @[Decoupled.scala 51:35]
  wire  _T_2 = axi_aw_ready & axi_aw_valid; // @[Decoupled.scala 51:35]
  wire  _T_3 = axi_w_ready & axi_w_valid; // @[Decoupled.scala 51:35]
  wire  _state_T = ~delay; // @[sram_AxiLite.scala 62:32]
  wire  _delay_T_1 = delay - 1'h1; // @[sram_AxiLite.scala 63:28]
  wire  _T_6 = 3'h2 == state; // @[sram_AxiLite.scala 47:20]
  wire  _state_T_2 = axi_r_ready & axi_r_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_3 = _state_T_2 ? 3'h0 : 3'h2; // @[sram_AxiLite.scala 66:25]
  wire [2:0] _state_T_5 = _state_T ? 3'h4 : 3'h3; // @[sram_AxiLite.scala 69:25]
  wire  _T_8 = 3'h4 == state; // @[sram_AxiLite.scala 47:20]
  wire  _state_T_6 = axi_b_ready & axi_b_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _state_T_7 = _state_T_6 ? 3'h0 : 3'h4; // @[sram_AxiLite.scala 73:25]
  wire [2:0] _GEN_2 = 3'h4 == state ? _state_T_7 : state; // @[sram_AxiLite.scala 47:20 73:19 46:24]
  wire [2:0] _GEN_3 = 3'h3 == state ? _state_T_5 : _GEN_2; // @[sram_AxiLite.scala 47:20 69:19]
  wire  _GEN_4 = 3'h3 == state ? _delay_T_1 : delay; // @[sram_AxiLite.scala 47:20 70:19 42:24]
  wire [31:0] _RamBB_i1_io_addr_T_1 = _T_6 ? axi_ar_bits_addr : 32'h0; // @[Mux.scala 81:58]
  RamBB RamBB_i1 ( // @[sram_AxiLite.scala 77:26]
    .clock(RamBB_i1_clock),
    .addr(RamBB_i1_addr),
    .mem_wen(RamBB_i1_mem_wen),
    .valid(RamBB_i1_valid),
    .wdata(RamBB_i1_wdata),
    .wmask(RamBB_i1_wmask),
    .rdata(RamBB_i1_rdata)
  );
  assign axi_ar_ready = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_r_valid = 3'h2 == state; // @[Mux.scala 81:61]
  assign axi_r_bits_data = RamBB_i1_rdata; // @[sram_AxiLite.scala 98:21]
  assign axi_aw_ready = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_w_ready = 3'h0 == state; // @[Mux.scala 81:61]
  assign axi_b_valid = 3'h4 == state; // @[Mux.scala 81:61]
  assign RamBB_i1_clock = clock; // @[sram_AxiLite.scala 78:25]
  assign RamBB_i1_addr = _T_8 ? axi_aw_bits_addr : _RamBB_i1_io_addr_T_1; // @[Mux.scala 81:58]
  assign RamBB_i1_mem_wen = 3'h4 == state; // @[Mux.scala 81:61]
  assign RamBB_i1_valid = _T_8 | _T_6; // @[Mux.scala 81:58]
  assign RamBB_i1_wdata = axi_w_bits_data; // @[sram_AxiLite.scala 92:25]
  assign RamBB_i1_wmask = axi_w_bits_strb; // @[sram_AxiLite.scala 93:25]
  always @(posedge clock) begin
    if (reset) begin // @[sram_AxiLite.scala 42:24]
      delay <= 1'h0; // @[sram_AxiLite.scala 42:24]
    end else if (3'h0 == state) begin // @[sram_AxiLite.scala 47:20]
      delay <= 1'h0; // @[sram_AxiLite.scala 49:19]
    end else if (3'h1 == state) begin // @[sram_AxiLite.scala 47:20]
      delay <= delay - 1'h1; // @[sram_AxiLite.scala 63:19]
    end else if (!(3'h2 == state)) begin // @[sram_AxiLite.scala 47:20]
      delay <= _GEN_4;
    end
    if (reset) begin // @[sram_AxiLite.scala 46:24]
      state <= 3'h0; // @[sram_AxiLite.scala 46:24]
    end else if (3'h0 == state) begin // @[sram_AxiLite.scala 47:20]
      if (_T_1) begin // @[sram_AxiLite.scala 51:32]
        state <= 3'h1; // @[sram_AxiLite.scala 52:23]
      end else if (_T_2 & _T_3) begin // @[sram_AxiLite.scala 54:51]
        state <= 3'h3; // @[sram_AxiLite.scala 55:23]
      end else begin
        state <= 3'h0; // @[sram_AxiLite.scala 58:23]
      end
    end else if (3'h1 == state) begin // @[sram_AxiLite.scala 47:20]
      if (~delay) begin // @[sram_AxiLite.scala 62:25]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[sram_AxiLite.scala 47:20]
      state <= _state_T_3; // @[sram_AxiLite.scala 66:19]
    end else begin
      state <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [31:0] io_out_inst,
  output [31:0] io_out_pc,
  output [31:0] io_out_difftest_mcause,
  output [31:0] io_out_difftest_mepc,
  output [31:0] io_out_difftest_mstatus,
  output [31:0] io_out_difftest_mtvec,
  output        io_out_wb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  IDU_i_from_IFU_valid; // @[core.scala 32:27]
  wire [31:0] IDU_i_from_IFU_bits_inst; // @[core.scala 32:27]
  wire [31:0] IDU_i_from_IFU_bits_pc; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_valid; // @[core.scala 32:27]
  wire [31:0] IDU_i_to_ISU_bits_imm; // @[core.scala 32:27]
  wire [31:0] IDU_i_to_ISU_bits_pc; // @[core.scala 32:27]
  wire [4:0] IDU_i_to_ISU_bits_rs1; // @[core.scala 32:27]
  wire [4:0] IDU_i_to_ISU_bits_rs2; // @[core.scala 32:27]
  wire [4:0] IDU_i_to_ISU_bits_rd; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_reg_wen; // @[core.scala 32:27]
  wire [2:0] IDU_i_to_ISU_bits_ctrl_sig_fu_op; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_mem_wen; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_is_ebreak; // @[core.scala 32:27]
  wire  IDU_i_to_ISU_bits_ctrl_sig_not_impl; // @[core.scala 32:27]
  wire [1:0] IDU_i_to_ISU_bits_ctrl_sig_src1_op; // @[core.scala 32:27]
  wire [1:0] IDU_i_to_ISU_bits_ctrl_sig_src2_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_alu_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_lsu_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_bru_op; // @[core.scala 32:27]
  wire [2:0] IDU_i_to_ISU_bits_ctrl_sig_csr_op; // @[core.scala 32:27]
  wire [3:0] IDU_i_to_ISU_bits_ctrl_sig_mdu_op; // @[core.scala 32:27]
  wire  ISU_i_clock; // @[core.scala 33:27]
  wire  ISU_i_reset; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_valid; // @[core.scala 33:27]
  wire [31:0] ISU_i_from_IDU_bits_imm; // @[core.scala 33:27]
  wire [31:0] ISU_i_from_IDU_bits_pc; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_IDU_bits_rs1; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_IDU_bits_rs2; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_IDU_bits_rd; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_reg_wen; // @[core.scala 33:27]
  wire [2:0] ISU_i_from_IDU_bits_ctrl_sig_fu_op; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_mem_wen; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_is_ebreak; // @[core.scala 33:27]
  wire  ISU_i_from_IDU_bits_ctrl_sig_not_impl; // @[core.scala 33:27]
  wire [1:0] ISU_i_from_IDU_bits_ctrl_sig_src1_op; // @[core.scala 33:27]
  wire [1:0] ISU_i_from_IDU_bits_ctrl_sig_src2_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_alu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_lsu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_bru_op; // @[core.scala 33:27]
  wire [2:0] ISU_i_from_IDU_bits_ctrl_sig_csr_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_from_IDU_bits_ctrl_sig_mdu_op; // @[core.scala 33:27]
  wire  ISU_i_from_WBU_bits_reg_wen; // @[core.scala 33:27]
  wire [31:0] ISU_i_from_WBU_bits_wdata; // @[core.scala 33:27]
  wire [4:0] ISU_i_from_WBU_bits_rd; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_valid; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_imm; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_pc; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_rdata1; // @[core.scala 33:27]
  wire [31:0] ISU_i_to_EXU_bits_rdata2; // @[core.scala 33:27]
  wire [4:0] ISU_i_to_EXU_bits_rd; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_reg_wen; // @[core.scala 33:27]
  wire [2:0] ISU_i_to_EXU_bits_ctrl_sig_fu_op; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_mem_wen; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_is_ebreak; // @[core.scala 33:27]
  wire  ISU_i_to_EXU_bits_ctrl_sig_not_impl; // @[core.scala 33:27]
  wire [1:0] ISU_i_to_EXU_bits_ctrl_sig_src1_op; // @[core.scala 33:27]
  wire [1:0] ISU_i_to_EXU_bits_ctrl_sig_src2_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_alu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_lsu_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_bru_op; // @[core.scala 33:27]
  wire [2:0] ISU_i_to_EXU_bits_ctrl_sig_csr_op; // @[core.scala 33:27]
  wire [3:0] ISU_i_to_EXU_bits_ctrl_sig_mdu_op; // @[core.scala 33:27]
  wire  EXU_i_clock; // @[core.scala 34:27]
  wire  EXU_i_reset; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_ready; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_imm; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_pc; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_rdata1; // @[core.scala 34:27]
  wire [31:0] EXU_i_from_ISU_bits_rdata2; // @[core.scala 34:27]
  wire [4:0] EXU_i_from_ISU_bits_rd; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_reg_wen; // @[core.scala 34:27]
  wire [2:0] EXU_i_from_ISU_bits_ctrl_sig_fu_op; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_mem_wen; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_is_ebreak; // @[core.scala 34:27]
  wire  EXU_i_from_ISU_bits_ctrl_sig_not_impl; // @[core.scala 34:27]
  wire [1:0] EXU_i_from_ISU_bits_ctrl_sig_src1_op; // @[core.scala 34:27]
  wire [1:0] EXU_i_from_ISU_bits_ctrl_sig_src2_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_alu_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_lsu_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_bru_op; // @[core.scala 34:27]
  wire [2:0] EXU_i_from_ISU_bits_ctrl_sig_csr_op; // @[core.scala 34:27]
  wire [3:0] EXU_i_from_ISU_bits_ctrl_sig_mdu_op; // @[core.scala 34:27]
  wire  EXU_i_to_WBU_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_alu_result; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_mdu_result; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_lsu_rdata; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_csr_rdata; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_WBU_bits_pc; // @[core.scala 34:27]
  wire  EXU_i_to_WBU_bits_reg_wen; // @[core.scala 34:27]
  wire [4:0] EXU_i_to_WBU_bits_rd; // @[core.scala 34:27]
  wire [2:0] EXU_i_to_WBU_bits_fu_op; // @[core.scala 34:27]
  wire  EXU_i_to_IFU_bits_bru_ctrl_br; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_IFU_bits_bru_addr; // @[core.scala 34:27]
  wire  EXU_i_to_IFU_bits_csr_ctrl_br; // @[core.scala 34:27]
  wire [31:0] EXU_i_to_IFU_bits_csr_addr; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mcause; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mepc; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mstatus; // @[core.scala 34:27]
  wire [31:0] EXU_i_difftest_mtvec; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_ar_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_ar_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_ar_bits_addr; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_r_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_r_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_r_bits_data; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_aw_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_aw_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_aw_bits_addr; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_w_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_w_valid; // @[core.scala 34:27]
  wire [31:0] EXU_i_lsu_axi_master_w_bits_data; // @[core.scala 34:27]
  wire [3:0] EXU_i_lsu_axi_master_w_bits_strb; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_b_ready; // @[core.scala 34:27]
  wire  EXU_i_lsu_axi_master_b_valid; // @[core.scala 34:27]
  wire  WBU_i_from_EXU_ready; // @[core.scala 35:27]
  wire  WBU_i_from_EXU_valid; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_alu_result; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_mdu_result; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_lsu_rdata; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_csr_rdata; // @[core.scala 35:27]
  wire [31:0] WBU_i_from_EXU_bits_pc; // @[core.scala 35:27]
  wire  WBU_i_from_EXU_bits_reg_wen; // @[core.scala 35:27]
  wire [4:0] WBU_i_from_EXU_bits_rd; // @[core.scala 35:27]
  wire [2:0] WBU_i_from_EXU_bits_fu_op; // @[core.scala 35:27]
  wire  WBU_i_to_ISU_bits_reg_wen; // @[core.scala 35:27]
  wire [31:0] WBU_i_to_ISU_bits_wdata; // @[core.scala 35:27]
  wire [4:0] WBU_i_to_ISU_bits_rd; // @[core.scala 35:27]
  wire  WBU_i_to_IFU_valid; // @[core.scala 35:27]
  wire  IFU_i_clock; // @[core.scala 48:27]
  wire  IFU_i_reset; // @[core.scala 48:27]
  wire  IFU_i_to_IDU_valid; // @[core.scala 48:27]
  wire [31:0] IFU_i_to_IDU_bits_inst; // @[core.scala 48:27]
  wire [31:0] IFU_i_to_IDU_bits_pc; // @[core.scala 48:27]
  wire  IFU_i_from_EXU_bits_bru_ctrl_br; // @[core.scala 48:27]
  wire [31:0] IFU_i_from_EXU_bits_bru_addr; // @[core.scala 48:27]
  wire  IFU_i_from_EXU_bits_csr_ctrl_br; // @[core.scala 48:27]
  wire [31:0] IFU_i_from_EXU_bits_csr_addr; // @[core.scala 48:27]
  wire  IFU_i_from_WBU_ready; // @[core.scala 48:27]
  wire  IFU_i_from_WBU_valid; // @[core.scala 48:27]
  wire  IFU_i_to_cache_ready; // @[core.scala 48:27]
  wire  IFU_i_to_cache_valid; // @[core.scala 48:27]
  wire [31:0] IFU_i_to_cache_bits_addr; // @[core.scala 48:27]
  wire  IFU_i_from_cache_ready; // @[core.scala 48:27]
  wire  IFU_i_from_cache_valid; // @[core.scala 48:27]
  wire [31:0] IFU_i_from_cache_bits_data; // @[core.scala 48:27]
  wire  icache_clock; // @[core.scala 49:27]
  wire  icache_reset; // @[core.scala 49:27]
  wire  icache_from_IFU_ready; // @[core.scala 49:27]
  wire  icache_from_IFU_valid; // @[core.scala 49:27]
  wire [31:0] icache_from_IFU_bits_addr; // @[core.scala 49:27]
  wire  icache_to_IFU_valid; // @[core.scala 49:27]
  wire [31:0] icache_to_IFU_bits_data; // @[core.scala 49:27]
  wire  icache_to_sram_ar_ready; // @[core.scala 49:27]
  wire  icache_to_sram_ar_valid; // @[core.scala 49:27]
  wire [31:0] icache_to_sram_ar_bits_addr; // @[core.scala 49:27]
  wire [7:0] icache_to_sram_ar_bits_len; // @[core.scala 49:27]
  wire  icache_to_sram_r_ready; // @[core.scala 49:27]
  wire  icache_to_sram_r_valid; // @[core.scala 49:27]
  wire [31:0] icache_to_sram_r_bits_data; // @[core.scala 49:27]
  wire  icache_to_sram_r_bits_last; // @[core.scala 49:27]
  wire  sram_i_clock; // @[core.scala 50:27]
  wire  sram_i_reset; // @[core.scala 50:27]
  wire  sram_i_axi_ar_ready; // @[core.scala 50:27]
  wire  sram_i_axi_ar_valid; // @[core.scala 50:27]
  wire [31:0] sram_i_axi_ar_bits_addr; // @[core.scala 50:27]
  wire [7:0] sram_i_axi_ar_bits_len; // @[core.scala 50:27]
  wire  sram_i_axi_r_ready; // @[core.scala 50:27]
  wire  sram_i_axi_r_valid; // @[core.scala 50:27]
  wire [31:0] sram_i_axi_r_bits_data; // @[core.scala 50:27]
  wire  sram_i_axi_r_bits_last; // @[core.scala 50:27]
  wire  sram_i2_clock; // @[core.scala 57:27]
  wire  sram_i2_reset; // @[core.scala 57:27]
  wire  sram_i2_axi_ar_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_ar_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_ar_bits_addr; // @[core.scala 57:27]
  wire  sram_i2_axi_r_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_r_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_r_bits_data; // @[core.scala 57:27]
  wire  sram_i2_axi_aw_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_aw_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_aw_bits_addr; // @[core.scala 57:27]
  wire  sram_i2_axi_w_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_w_valid; // @[core.scala 57:27]
  wire [31:0] sram_i2_axi_w_bits_data; // @[core.scala 57:27]
  wire [3:0] sram_i2_axi_w_bits_strb; // @[core.scala 57:27]
  wire  sram_i2_axi_b_ready; // @[core.scala 57:27]
  wire  sram_i2_axi_b_valid; // @[core.scala 57:27]
  wire  _EXU_i_from_ISU_bits_T = ISU_i_to_EXU_valid & EXU_i_from_ISU_ready; // @[Connect.scala 26:58]
  reg [31:0] EXU_i_from_ISU_bits_r_imm; // @[Reg.scala 19:16]
  reg [31:0] EXU_i_from_ISU_bits_r_pc; // @[Reg.scala 19:16]
  reg [31:0] EXU_i_from_ISU_bits_r_rdata1; // @[Reg.scala 19:16]
  reg [31:0] EXU_i_from_ISU_bits_r_rdata2; // @[Reg.scala 19:16]
  reg [4:0] EXU_i_from_ISU_bits_r_rd; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen; // @[Reg.scala 19:16]
  reg [2:0] EXU_i_from_ISU_bits_r_ctrl_sig_fu_op; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak; // @[Reg.scala 19:16]
  reg  EXU_i_from_ISU_bits_r_ctrl_sig_not_impl; // @[Reg.scala 19:16]
  reg [1:0] EXU_i_from_ISU_bits_r_ctrl_sig_src1_op; // @[Reg.scala 19:16]
  reg [1:0] EXU_i_from_ISU_bits_r_ctrl_sig_src2_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_alu_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_bru_op; // @[Reg.scala 19:16]
  reg [2:0] EXU_i_from_ISU_bits_r_ctrl_sig_csr_op; // @[Reg.scala 19:16]
  reg [3:0] EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op; // @[Reg.scala 19:16]
  IDU IDU_i ( // @[core.scala 32:27]
    .from_IFU_valid(IDU_i_from_IFU_valid),
    .from_IFU_bits_inst(IDU_i_from_IFU_bits_inst),
    .from_IFU_bits_pc(IDU_i_from_IFU_bits_pc),
    .to_ISU_valid(IDU_i_to_ISU_valid),
    .to_ISU_bits_imm(IDU_i_to_ISU_bits_imm),
    .to_ISU_bits_pc(IDU_i_to_ISU_bits_pc),
    .to_ISU_bits_rs1(IDU_i_to_ISU_bits_rs1),
    .to_ISU_bits_rs2(IDU_i_to_ISU_bits_rs2),
    .to_ISU_bits_rd(IDU_i_to_ISU_bits_rd),
    .to_ISU_bits_ctrl_sig_reg_wen(IDU_i_to_ISU_bits_ctrl_sig_reg_wen),
    .to_ISU_bits_ctrl_sig_fu_op(IDU_i_to_ISU_bits_ctrl_sig_fu_op),
    .to_ISU_bits_ctrl_sig_mem_wen(IDU_i_to_ISU_bits_ctrl_sig_mem_wen),
    .to_ISU_bits_ctrl_sig_is_ebreak(IDU_i_to_ISU_bits_ctrl_sig_is_ebreak),
    .to_ISU_bits_ctrl_sig_not_impl(IDU_i_to_ISU_bits_ctrl_sig_not_impl),
    .to_ISU_bits_ctrl_sig_src1_op(IDU_i_to_ISU_bits_ctrl_sig_src1_op),
    .to_ISU_bits_ctrl_sig_src2_op(IDU_i_to_ISU_bits_ctrl_sig_src2_op),
    .to_ISU_bits_ctrl_sig_alu_op(IDU_i_to_ISU_bits_ctrl_sig_alu_op),
    .to_ISU_bits_ctrl_sig_lsu_op(IDU_i_to_ISU_bits_ctrl_sig_lsu_op),
    .to_ISU_bits_ctrl_sig_bru_op(IDU_i_to_ISU_bits_ctrl_sig_bru_op),
    .to_ISU_bits_ctrl_sig_csr_op(IDU_i_to_ISU_bits_ctrl_sig_csr_op),
    .to_ISU_bits_ctrl_sig_mdu_op(IDU_i_to_ISU_bits_ctrl_sig_mdu_op)
  );
  ISU ISU_i ( // @[core.scala 33:27]
    .clock(ISU_i_clock),
    .reset(ISU_i_reset),
    .from_IDU_valid(ISU_i_from_IDU_valid),
    .from_IDU_bits_imm(ISU_i_from_IDU_bits_imm),
    .from_IDU_bits_pc(ISU_i_from_IDU_bits_pc),
    .from_IDU_bits_rs1(ISU_i_from_IDU_bits_rs1),
    .from_IDU_bits_rs2(ISU_i_from_IDU_bits_rs2),
    .from_IDU_bits_rd(ISU_i_from_IDU_bits_rd),
    .from_IDU_bits_ctrl_sig_reg_wen(ISU_i_from_IDU_bits_ctrl_sig_reg_wen),
    .from_IDU_bits_ctrl_sig_fu_op(ISU_i_from_IDU_bits_ctrl_sig_fu_op),
    .from_IDU_bits_ctrl_sig_mem_wen(ISU_i_from_IDU_bits_ctrl_sig_mem_wen),
    .from_IDU_bits_ctrl_sig_is_ebreak(ISU_i_from_IDU_bits_ctrl_sig_is_ebreak),
    .from_IDU_bits_ctrl_sig_not_impl(ISU_i_from_IDU_bits_ctrl_sig_not_impl),
    .from_IDU_bits_ctrl_sig_src1_op(ISU_i_from_IDU_bits_ctrl_sig_src1_op),
    .from_IDU_bits_ctrl_sig_src2_op(ISU_i_from_IDU_bits_ctrl_sig_src2_op),
    .from_IDU_bits_ctrl_sig_alu_op(ISU_i_from_IDU_bits_ctrl_sig_alu_op),
    .from_IDU_bits_ctrl_sig_lsu_op(ISU_i_from_IDU_bits_ctrl_sig_lsu_op),
    .from_IDU_bits_ctrl_sig_bru_op(ISU_i_from_IDU_bits_ctrl_sig_bru_op),
    .from_IDU_bits_ctrl_sig_csr_op(ISU_i_from_IDU_bits_ctrl_sig_csr_op),
    .from_IDU_bits_ctrl_sig_mdu_op(ISU_i_from_IDU_bits_ctrl_sig_mdu_op),
    .from_WBU_bits_reg_wen(ISU_i_from_WBU_bits_reg_wen),
    .from_WBU_bits_wdata(ISU_i_from_WBU_bits_wdata),
    .from_WBU_bits_rd(ISU_i_from_WBU_bits_rd),
    .to_EXU_valid(ISU_i_to_EXU_valid),
    .to_EXU_bits_imm(ISU_i_to_EXU_bits_imm),
    .to_EXU_bits_pc(ISU_i_to_EXU_bits_pc),
    .to_EXU_bits_rdata1(ISU_i_to_EXU_bits_rdata1),
    .to_EXU_bits_rdata2(ISU_i_to_EXU_bits_rdata2),
    .to_EXU_bits_rd(ISU_i_to_EXU_bits_rd),
    .to_EXU_bits_ctrl_sig_reg_wen(ISU_i_to_EXU_bits_ctrl_sig_reg_wen),
    .to_EXU_bits_ctrl_sig_fu_op(ISU_i_to_EXU_bits_ctrl_sig_fu_op),
    .to_EXU_bits_ctrl_sig_mem_wen(ISU_i_to_EXU_bits_ctrl_sig_mem_wen),
    .to_EXU_bits_ctrl_sig_is_ebreak(ISU_i_to_EXU_bits_ctrl_sig_is_ebreak),
    .to_EXU_bits_ctrl_sig_not_impl(ISU_i_to_EXU_bits_ctrl_sig_not_impl),
    .to_EXU_bits_ctrl_sig_src1_op(ISU_i_to_EXU_bits_ctrl_sig_src1_op),
    .to_EXU_bits_ctrl_sig_src2_op(ISU_i_to_EXU_bits_ctrl_sig_src2_op),
    .to_EXU_bits_ctrl_sig_alu_op(ISU_i_to_EXU_bits_ctrl_sig_alu_op),
    .to_EXU_bits_ctrl_sig_lsu_op(ISU_i_to_EXU_bits_ctrl_sig_lsu_op),
    .to_EXU_bits_ctrl_sig_bru_op(ISU_i_to_EXU_bits_ctrl_sig_bru_op),
    .to_EXU_bits_ctrl_sig_csr_op(ISU_i_to_EXU_bits_ctrl_sig_csr_op),
    .to_EXU_bits_ctrl_sig_mdu_op(ISU_i_to_EXU_bits_ctrl_sig_mdu_op)
  );
  EXU EXU_i ( // @[core.scala 34:27]
    .clock(EXU_i_clock),
    .reset(EXU_i_reset),
    .from_ISU_ready(EXU_i_from_ISU_ready),
    .from_ISU_valid(EXU_i_from_ISU_valid),
    .from_ISU_bits_imm(EXU_i_from_ISU_bits_imm),
    .from_ISU_bits_pc(EXU_i_from_ISU_bits_pc),
    .from_ISU_bits_rdata1(EXU_i_from_ISU_bits_rdata1),
    .from_ISU_bits_rdata2(EXU_i_from_ISU_bits_rdata2),
    .from_ISU_bits_rd(EXU_i_from_ISU_bits_rd),
    .from_ISU_bits_ctrl_sig_reg_wen(EXU_i_from_ISU_bits_ctrl_sig_reg_wen),
    .from_ISU_bits_ctrl_sig_fu_op(EXU_i_from_ISU_bits_ctrl_sig_fu_op),
    .from_ISU_bits_ctrl_sig_mem_wen(EXU_i_from_ISU_bits_ctrl_sig_mem_wen),
    .from_ISU_bits_ctrl_sig_is_ebreak(EXU_i_from_ISU_bits_ctrl_sig_is_ebreak),
    .from_ISU_bits_ctrl_sig_not_impl(EXU_i_from_ISU_bits_ctrl_sig_not_impl),
    .from_ISU_bits_ctrl_sig_src1_op(EXU_i_from_ISU_bits_ctrl_sig_src1_op),
    .from_ISU_bits_ctrl_sig_src2_op(EXU_i_from_ISU_bits_ctrl_sig_src2_op),
    .from_ISU_bits_ctrl_sig_alu_op(EXU_i_from_ISU_bits_ctrl_sig_alu_op),
    .from_ISU_bits_ctrl_sig_lsu_op(EXU_i_from_ISU_bits_ctrl_sig_lsu_op),
    .from_ISU_bits_ctrl_sig_bru_op(EXU_i_from_ISU_bits_ctrl_sig_bru_op),
    .from_ISU_bits_ctrl_sig_csr_op(EXU_i_from_ISU_bits_ctrl_sig_csr_op),
    .from_ISU_bits_ctrl_sig_mdu_op(EXU_i_from_ISU_bits_ctrl_sig_mdu_op),
    .to_WBU_valid(EXU_i_to_WBU_valid),
    .to_WBU_bits_alu_result(EXU_i_to_WBU_bits_alu_result),
    .to_WBU_bits_mdu_result(EXU_i_to_WBU_bits_mdu_result),
    .to_WBU_bits_lsu_rdata(EXU_i_to_WBU_bits_lsu_rdata),
    .to_WBU_bits_csr_rdata(EXU_i_to_WBU_bits_csr_rdata),
    .to_WBU_bits_pc(EXU_i_to_WBU_bits_pc),
    .to_WBU_bits_reg_wen(EXU_i_to_WBU_bits_reg_wen),
    .to_WBU_bits_rd(EXU_i_to_WBU_bits_rd),
    .to_WBU_bits_fu_op(EXU_i_to_WBU_bits_fu_op),
    .to_IFU_bits_bru_ctrl_br(EXU_i_to_IFU_bits_bru_ctrl_br),
    .to_IFU_bits_bru_addr(EXU_i_to_IFU_bits_bru_addr),
    .to_IFU_bits_csr_ctrl_br(EXU_i_to_IFU_bits_csr_ctrl_br),
    .to_IFU_bits_csr_addr(EXU_i_to_IFU_bits_csr_addr),
    .difftest_mcause(EXU_i_difftest_mcause),
    .difftest_mepc(EXU_i_difftest_mepc),
    .difftest_mstatus(EXU_i_difftest_mstatus),
    .difftest_mtvec(EXU_i_difftest_mtvec),
    .lsu_axi_master_ar_ready(EXU_i_lsu_axi_master_ar_ready),
    .lsu_axi_master_ar_valid(EXU_i_lsu_axi_master_ar_valid),
    .lsu_axi_master_ar_bits_addr(EXU_i_lsu_axi_master_ar_bits_addr),
    .lsu_axi_master_r_ready(EXU_i_lsu_axi_master_r_ready),
    .lsu_axi_master_r_valid(EXU_i_lsu_axi_master_r_valid),
    .lsu_axi_master_r_bits_data(EXU_i_lsu_axi_master_r_bits_data),
    .lsu_axi_master_aw_ready(EXU_i_lsu_axi_master_aw_ready),
    .lsu_axi_master_aw_valid(EXU_i_lsu_axi_master_aw_valid),
    .lsu_axi_master_aw_bits_addr(EXU_i_lsu_axi_master_aw_bits_addr),
    .lsu_axi_master_w_ready(EXU_i_lsu_axi_master_w_ready),
    .lsu_axi_master_w_valid(EXU_i_lsu_axi_master_w_valid),
    .lsu_axi_master_w_bits_data(EXU_i_lsu_axi_master_w_bits_data),
    .lsu_axi_master_w_bits_strb(EXU_i_lsu_axi_master_w_bits_strb),
    .lsu_axi_master_b_ready(EXU_i_lsu_axi_master_b_ready),
    .lsu_axi_master_b_valid(EXU_i_lsu_axi_master_b_valid)
  );
  WBU WBU_i ( // @[core.scala 35:27]
    .from_EXU_ready(WBU_i_from_EXU_ready),
    .from_EXU_valid(WBU_i_from_EXU_valid),
    .from_EXU_bits_alu_result(WBU_i_from_EXU_bits_alu_result),
    .from_EXU_bits_mdu_result(WBU_i_from_EXU_bits_mdu_result),
    .from_EXU_bits_lsu_rdata(WBU_i_from_EXU_bits_lsu_rdata),
    .from_EXU_bits_csr_rdata(WBU_i_from_EXU_bits_csr_rdata),
    .from_EXU_bits_pc(WBU_i_from_EXU_bits_pc),
    .from_EXU_bits_reg_wen(WBU_i_from_EXU_bits_reg_wen),
    .from_EXU_bits_rd(WBU_i_from_EXU_bits_rd),
    .from_EXU_bits_fu_op(WBU_i_from_EXU_bits_fu_op),
    .to_ISU_bits_reg_wen(WBU_i_to_ISU_bits_reg_wen),
    .to_ISU_bits_wdata(WBU_i_to_ISU_bits_wdata),
    .to_ISU_bits_rd(WBU_i_to_ISU_bits_rd),
    .to_IFU_valid(WBU_i_to_IFU_valid)
  );
  IFU_cache IFU_i ( // @[core.scala 48:27]
    .clock(IFU_i_clock),
    .reset(IFU_i_reset),
    .to_IDU_valid(IFU_i_to_IDU_valid),
    .to_IDU_bits_inst(IFU_i_to_IDU_bits_inst),
    .to_IDU_bits_pc(IFU_i_to_IDU_bits_pc),
    .from_EXU_bits_bru_ctrl_br(IFU_i_from_EXU_bits_bru_ctrl_br),
    .from_EXU_bits_bru_addr(IFU_i_from_EXU_bits_bru_addr),
    .from_EXU_bits_csr_ctrl_br(IFU_i_from_EXU_bits_csr_ctrl_br),
    .from_EXU_bits_csr_addr(IFU_i_from_EXU_bits_csr_addr),
    .from_WBU_ready(IFU_i_from_WBU_ready),
    .from_WBU_valid(IFU_i_from_WBU_valid),
    .to_cache_ready(IFU_i_to_cache_ready),
    .to_cache_valid(IFU_i_to_cache_valid),
    .to_cache_bits_addr(IFU_i_to_cache_bits_addr),
    .from_cache_ready(IFU_i_from_cache_ready),
    .from_cache_valid(IFU_i_from_cache_valid),
    .from_cache_bits_data(IFU_i_from_cache_bits_data)
  );
  I_Cache icache ( // @[core.scala 49:27]
    .clock(icache_clock),
    .reset(icache_reset),
    .from_IFU_ready(icache_from_IFU_ready),
    .from_IFU_valid(icache_from_IFU_valid),
    .from_IFU_bits_addr(icache_from_IFU_bits_addr),
    .to_IFU_valid(icache_to_IFU_valid),
    .to_IFU_bits_data(icache_to_IFU_bits_data),
    .to_sram_ar_ready(icache_to_sram_ar_ready),
    .to_sram_ar_valid(icache_to_sram_ar_valid),
    .to_sram_ar_bits_addr(icache_to_sram_ar_bits_addr),
    .to_sram_ar_bits_len(icache_to_sram_ar_bits_len),
    .to_sram_r_ready(icache_to_sram_r_ready),
    .to_sram_r_valid(icache_to_sram_r_valid),
    .to_sram_r_bits_data(icache_to_sram_r_bits_data),
    .to_sram_r_bits_last(icache_to_sram_r_bits_last)
  );
  SRAM_axi sram_i ( // @[core.scala 50:27]
    .clock(sram_i_clock),
    .reset(sram_i_reset),
    .axi_ar_ready(sram_i_axi_ar_ready),
    .axi_ar_valid(sram_i_axi_ar_valid),
    .axi_ar_bits_addr(sram_i_axi_ar_bits_addr),
    .axi_ar_bits_len(sram_i_axi_ar_bits_len),
    .axi_r_ready(sram_i_axi_r_ready),
    .axi_r_valid(sram_i_axi_r_valid),
    .axi_r_bits_data(sram_i_axi_r_bits_data),
    .axi_r_bits_last(sram_i_axi_r_bits_last)
  );
  SRAM sram_i2 ( // @[core.scala 57:27]
    .clock(sram_i2_clock),
    .reset(sram_i2_reset),
    .axi_ar_ready(sram_i2_axi_ar_ready),
    .axi_ar_valid(sram_i2_axi_ar_valid),
    .axi_ar_bits_addr(sram_i2_axi_ar_bits_addr),
    .axi_r_ready(sram_i2_axi_r_ready),
    .axi_r_valid(sram_i2_axi_r_valid),
    .axi_r_bits_data(sram_i2_axi_r_bits_data),
    .axi_aw_ready(sram_i2_axi_aw_ready),
    .axi_aw_valid(sram_i2_axi_aw_valid),
    .axi_aw_bits_addr(sram_i2_axi_aw_bits_addr),
    .axi_w_ready(sram_i2_axi_w_ready),
    .axi_w_valid(sram_i2_axi_w_valid),
    .axi_w_bits_data(sram_i2_axi_w_bits_data),
    .axi_w_bits_strb(sram_i2_axi_w_bits_strb),
    .axi_b_ready(sram_i2_axi_b_ready),
    .axi_b_valid(sram_i2_axi_b_valid)
  );
  assign io_out_inst = IFU_i_to_IDU_bits_inst; // @[core.scala 75:20]
  assign io_out_pc = IFU_i_to_IDU_bits_pc; // @[core.scala 76:20]
  assign io_out_difftest_mcause = EXU_i_difftest_mcause; // @[core.scala 79:21]
  assign io_out_difftest_mepc = EXU_i_difftest_mepc; // @[core.scala 79:21]
  assign io_out_difftest_mstatus = EXU_i_difftest_mstatus; // @[core.scala 79:21]
  assign io_out_difftest_mtvec = EXU_i_difftest_mtvec; // @[core.scala 79:21]
  assign io_out_wb = WBU_i_to_IFU_valid; // @[core.scala 77:20]
  assign IDU_i_from_IFU_valid = IFU_i_to_IDU_valid; // @[Connect.scala 16:22]
  assign IDU_i_from_IFU_bits_inst = IFU_i_to_IDU_bits_inst; // @[Connect.scala 15:22]
  assign IDU_i_from_IFU_bits_pc = IFU_i_to_IDU_bits_pc; // @[Connect.scala 15:22]
  assign ISU_i_clock = clock;
  assign ISU_i_reset = reset;
  assign ISU_i_from_IDU_valid = IDU_i_to_ISU_valid; // @[Connect.scala 16:22]
  assign ISU_i_from_IDU_bits_imm = IDU_i_to_ISU_bits_imm; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_pc = IDU_i_to_ISU_bits_pc; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_rs1 = IDU_i_to_ISU_bits_rs1; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_rs2 = IDU_i_to_ISU_bits_rs2; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_rd = IDU_i_to_ISU_bits_rd; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_reg_wen = IDU_i_to_ISU_bits_ctrl_sig_reg_wen; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_fu_op = IDU_i_to_ISU_bits_ctrl_sig_fu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_mem_wen = IDU_i_to_ISU_bits_ctrl_sig_mem_wen; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_is_ebreak = IDU_i_to_ISU_bits_ctrl_sig_is_ebreak; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_not_impl = IDU_i_to_ISU_bits_ctrl_sig_not_impl; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_src1_op = IDU_i_to_ISU_bits_ctrl_sig_src1_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_src2_op = IDU_i_to_ISU_bits_ctrl_sig_src2_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_alu_op = IDU_i_to_ISU_bits_ctrl_sig_alu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_lsu_op = IDU_i_to_ISU_bits_ctrl_sig_lsu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_bru_op = IDU_i_to_ISU_bits_ctrl_sig_bru_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_csr_op = IDU_i_to_ISU_bits_ctrl_sig_csr_op; // @[Connect.scala 15:22]
  assign ISU_i_from_IDU_bits_ctrl_sig_mdu_op = IDU_i_to_ISU_bits_ctrl_sig_mdu_op; // @[Connect.scala 15:22]
  assign ISU_i_from_WBU_bits_reg_wen = WBU_i_to_ISU_bits_reg_wen; // @[Connect.scala 15:22]
  assign ISU_i_from_WBU_bits_wdata = WBU_i_to_ISU_bits_wdata; // @[Connect.scala 15:22]
  assign ISU_i_from_WBU_bits_rd = WBU_i_to_ISU_bits_rd; // @[Connect.scala 15:22]
  assign EXU_i_clock = clock;
  assign EXU_i_reset = reset;
  assign EXU_i_from_ISU_valid = ISU_i_to_EXU_valid; // @[Connect.scala 27:22]
  assign EXU_i_from_ISU_bits_imm = EXU_i_from_ISU_bits_r_imm; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_pc = EXU_i_from_ISU_bits_r_pc; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_rdata1 = EXU_i_from_ISU_bits_r_rdata1; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_rdata2 = EXU_i_from_ISU_bits_r_rdata2; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_rd = EXU_i_from_ISU_bits_r_rd; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_reg_wen = EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_fu_op = EXU_i_from_ISU_bits_r_ctrl_sig_fu_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_mem_wen = EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_is_ebreak = EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_not_impl = EXU_i_from_ISU_bits_r_ctrl_sig_not_impl; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_src1_op = EXU_i_from_ISU_bits_r_ctrl_sig_src1_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_src2_op = EXU_i_from_ISU_bits_r_ctrl_sig_src2_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_alu_op = EXU_i_from_ISU_bits_r_ctrl_sig_alu_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_lsu_op = EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_bru_op = EXU_i_from_ISU_bits_r_ctrl_sig_bru_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_csr_op = EXU_i_from_ISU_bits_r_ctrl_sig_csr_op; // @[Connect.scala 26:22]
  assign EXU_i_from_ISU_bits_ctrl_sig_mdu_op = EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op; // @[Connect.scala 26:22]
  assign EXU_i_lsu_axi_master_ar_ready = sram_i2_axi_ar_ready; // @[Connect.scala 17:22]
  assign EXU_i_lsu_axi_master_r_valid = sram_i2_axi_r_valid; // @[Connect.scala 16:22]
  assign EXU_i_lsu_axi_master_r_bits_data = sram_i2_axi_r_bits_data; // @[Connect.scala 15:22]
  assign EXU_i_lsu_axi_master_aw_ready = sram_i2_axi_aw_ready; // @[Connect.scala 17:22]
  assign EXU_i_lsu_axi_master_w_ready = sram_i2_axi_w_ready; // @[Connect.scala 17:22]
  assign EXU_i_lsu_axi_master_b_valid = sram_i2_axi_b_valid; // @[Connect.scala 16:22]
  assign WBU_i_from_EXU_valid = EXU_i_to_WBU_valid; // @[Connect.scala 16:22]
  assign WBU_i_from_EXU_bits_alu_result = EXU_i_to_WBU_bits_alu_result; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_mdu_result = EXU_i_to_WBU_bits_mdu_result; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_lsu_rdata = EXU_i_to_WBU_bits_lsu_rdata; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_csr_rdata = EXU_i_to_WBU_bits_csr_rdata; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_pc = EXU_i_to_WBU_bits_pc; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_reg_wen = EXU_i_to_WBU_bits_reg_wen; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_rd = EXU_i_to_WBU_bits_rd; // @[Connect.scala 15:22]
  assign WBU_i_from_EXU_bits_fu_op = EXU_i_to_WBU_bits_fu_op; // @[Connect.scala 15:22]
  assign IFU_i_clock = clock;
  assign IFU_i_reset = reset;
  assign IFU_i_from_EXU_bits_bru_ctrl_br = EXU_i_to_IFU_bits_bru_ctrl_br; // @[Connect.scala 15:22]
  assign IFU_i_from_EXU_bits_bru_addr = EXU_i_to_IFU_bits_bru_addr; // @[Connect.scala 15:22]
  assign IFU_i_from_EXU_bits_csr_ctrl_br = EXU_i_to_IFU_bits_csr_ctrl_br; // @[Connect.scala 15:22]
  assign IFU_i_from_EXU_bits_csr_addr = EXU_i_to_IFU_bits_csr_addr; // @[Connect.scala 15:22]
  assign IFU_i_from_WBU_valid = WBU_i_to_IFU_valid; // @[Connect.scala 16:22]
  assign IFU_i_to_cache_ready = icache_from_IFU_ready; // @[Connect.scala 17:22]
  assign IFU_i_from_cache_valid = icache_to_IFU_valid; // @[Connect.scala 16:22]
  assign IFU_i_from_cache_bits_data = icache_to_IFU_bits_data; // @[Connect.scala 15:22]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_from_IFU_valid = IFU_i_to_cache_valid; // @[Connect.scala 16:22]
  assign icache_from_IFU_bits_addr = IFU_i_to_cache_bits_addr; // @[Connect.scala 15:22]
  assign icache_to_sram_ar_ready = sram_i_axi_ar_ready; // @[Connect.scala 17:22]
  assign icache_to_sram_r_valid = sram_i_axi_r_valid; // @[Connect.scala 16:22]
  assign icache_to_sram_r_bits_data = sram_i_axi_r_bits_data; // @[Connect.scala 15:22]
  assign icache_to_sram_r_bits_last = sram_i_axi_r_bits_last; // @[Connect.scala 15:22]
  assign sram_i_clock = clock;
  assign sram_i_reset = reset;
  assign sram_i_axi_ar_valid = icache_to_sram_ar_valid; // @[Connect.scala 16:22]
  assign sram_i_axi_ar_bits_addr = icache_to_sram_ar_bits_addr; // @[Connect.scala 15:22]
  assign sram_i_axi_ar_bits_len = icache_to_sram_ar_bits_len; // @[Connect.scala 15:22]
  assign sram_i_axi_r_ready = icache_to_sram_r_ready; // @[Connect.scala 17:22]
  assign sram_i2_clock = clock;
  assign sram_i2_reset = reset;
  assign sram_i2_axi_ar_valid = EXU_i_lsu_axi_master_ar_valid; // @[Connect.scala 16:22]
  assign sram_i2_axi_ar_bits_addr = EXU_i_lsu_axi_master_ar_bits_addr; // @[Connect.scala 15:22]
  assign sram_i2_axi_r_ready = EXU_i_lsu_axi_master_r_ready; // @[Connect.scala 17:22]
  assign sram_i2_axi_aw_valid = EXU_i_lsu_axi_master_aw_valid; // @[Connect.scala 16:22]
  assign sram_i2_axi_aw_bits_addr = EXU_i_lsu_axi_master_aw_bits_addr; // @[Connect.scala 15:22]
  assign sram_i2_axi_w_valid = EXU_i_lsu_axi_master_w_valid; // @[Connect.scala 16:22]
  assign sram_i2_axi_w_bits_data = EXU_i_lsu_axi_master_w_bits_data; // @[Connect.scala 15:22]
  assign sram_i2_axi_w_bits_strb = EXU_i_lsu_axi_master_w_bits_strb; // @[Connect.scala 15:22]
  assign sram_i2_axi_b_ready = EXU_i_lsu_axi_master_b_ready; // @[Connect.scala 17:22]
  always @(posedge clock) begin
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_imm <= ISU_i_to_EXU_bits_imm; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_pc <= ISU_i_to_EXU_bits_pc; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_rdata1 <= ISU_i_to_EXU_bits_rdata1; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_rdata2 <= ISU_i_to_EXU_bits_rdata2; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_rd <= ISU_i_to_EXU_bits_rd; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen <= ISU_i_to_EXU_bits_ctrl_sig_reg_wen; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_fu_op <= ISU_i_to_EXU_bits_ctrl_sig_fu_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen <= ISU_i_to_EXU_bits_ctrl_sig_mem_wen; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak <= ISU_i_to_EXU_bits_ctrl_sig_is_ebreak; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_not_impl <= ISU_i_to_EXU_bits_ctrl_sig_not_impl; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_src1_op <= ISU_i_to_EXU_bits_ctrl_sig_src1_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_src2_op <= ISU_i_to_EXU_bits_ctrl_sig_src2_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_alu_op <= ISU_i_to_EXU_bits_ctrl_sig_alu_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op <= ISU_i_to_EXU_bits_ctrl_sig_lsu_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_bru_op <= ISU_i_to_EXU_bits_ctrl_sig_bru_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_csr_op <= ISU_i_to_EXU_bits_ctrl_sig_csr_op; // @[Reg.scala 20:22]
    end
    if (_EXU_i_from_ISU_bits_T) begin // @[Reg.scala 20:18]
      EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op <= ISU_i_to_EXU_bits_ctrl_sig_mdu_op; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_imm = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_rdata1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_rdata2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_rd = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_reg_wen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_fu_op = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_mem_wen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_is_ebreak = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_not_impl = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_src1_op = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_src2_op = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_alu_op = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_lsu_op = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_bru_op = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_csr_op = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  EXU_i_from_ISU_bits_r_ctrl_sig_mdu_op = _RAND_16[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
